magic
tech gf180mcuD
magscale 1 10
timestamp 1756715696
<< nwell >>
rect 1232 -119 1478 253
rect 1483 -119 1535 253
rect 2579 -119 2823 253
rect 1181 -239 1552 -119
rect 2512 -239 2883 -119
rect 1232 -266 1478 -239
rect 1483 -265 1535 -239
rect 2579 -265 2823 -239
<< pwell >>
rect 995 454 1051 971
rect 1273 673 1519 772
rect 2583 675 2827 771
rect 2513 673 2927 675
rect 1273 665 1582 673
rect 1186 545 1582 665
rect 2513 545 2941 673
rect 1273 465 1582 545
rect 1145 454 1582 465
rect 995 409 1582 454
rect 1012 348 1158 409
rect 1273 364 1582 409
rect 1273 348 1519 364
rect 1012 293 1519 348
rect 1012 254 1158 293
rect 1273 253 1582 293
rect 2583 253 2827 545
rect 2854 253 2941 545
rect 3585 253 4835 547
<< nsubdiff >>
rect 84 1533 184 1559
rect 84 1477 103 1533
rect 159 1477 184 1533
rect 84 1459 184 1477
rect 3434 -151 3534 -128
rect 3434 -207 3456 -151
rect 3512 -207 3534 -151
rect 3434 -228 3534 -207
<< nsubdiffcont >>
rect 103 1477 159 1533
rect 3456 -207 3512 -151
<< metal1 >>
rect 204 1079 392 1155
rect 3973 1053 4029 1472
rect 4455 1053 4511 1411
rect 3963 977 4039 1053
rect 4445 977 4521 1053
rect 3052 909 3193 929
rect 3052 853 3064 909
rect 3120 853 3193 909
rect 3052 835 3193 853
rect 3996 893 4488 903
rect 3996 837 4423 893
rect 4479 837 4488 893
rect 3996 827 4488 837
rect 1186 643 1259 665
rect 1483 665 1525 678
rect 2854 675 2901 685
rect 1320 643 1525 665
rect 1186 545 1525 643
rect 2513 545 2927 675
rect 3533 545 3745 665
rect 206 149 278 402
rect 779 348 822 357
rect 1661 348 1788 357
rect 430 -73 502 319
rect 779 293 1788 348
rect 1638 181 2320 245
rect 1181 -239 1552 -119
rect 2512 -153 2892 -119
rect 2512 -209 2661 -153
rect 2717 -209 2892 -153
rect 2512 -239 2892 -209
<< via1 >>
rect 2660 1484 2716 1540
rect 3291 1134 3347 1190
rect 4138 1134 4194 1190
rect 4290 1134 4346 1190
rect 995 985 1051 1041
rect 3064 853 3120 909
rect 4423 837 4479 893
rect 1259 643 1320 703
rect 1966 409 2022 465
rect 3023 195 3079 251
rect 3352 193 3408 249
rect 2661 -209 2717 -153
<< metal2 >>
rect 2638 1540 2731 1556
rect 2638 1484 2660 1540
rect 2716 1484 2731 1540
rect 2638 1468 2731 1484
rect 3280 1190 3356 1200
rect 4128 1190 4204 1199
rect 3280 1134 3291 1190
rect 3347 1134 4138 1190
rect 4194 1134 4204 1190
rect 3280 1124 3356 1134
rect 4128 1123 4204 1134
rect 4280 1190 4356 1199
rect 4280 1134 4290 1190
rect 4346 1134 4356 1190
rect 4280 1123 4356 1134
rect 984 1041 1060 1050
rect 984 985 995 1041
rect 1051 985 1060 1041
rect 984 974 1060 985
rect 995 465 1051 974
rect 3023 909 3132 921
rect 3023 853 3064 909
rect 3120 853 3132 909
rect 3023 841 3132 853
rect 1232 703 1344 728
rect 1232 643 1259 703
rect 1320 643 1344 703
rect 1232 616 1344 643
rect 1957 465 2033 477
rect 995 409 1966 465
rect 2022 409 2033 465
rect 1957 401 2033 409
rect 3023 263 3079 841
rect 3011 251 3091 263
rect 3011 195 3023 251
rect 3079 195 3091 251
rect 3011 186 3091 195
rect 3342 249 3418 261
rect 4290 249 4346 1123
rect 4412 893 4488 903
rect 4412 837 4423 893
rect 4479 837 4488 893
rect 4412 827 4488 837
rect 3342 193 3352 249
rect 3408 193 4346 249
rect 3342 185 3418 193
rect 4423 -53 4479 827
rect 2649 -153 2725 -142
rect 2649 -209 2661 -153
rect 2717 -209 2725 -153
rect 2649 -218 2725 -209
<< via2 >>
rect 2660 1484 2716 1540
rect 1259 643 1320 703
rect 2661 -209 2717 -153
<< metal3 >>
rect 1176 703 1400 2603
rect 1176 643 1259 703
rect 1320 643 1400 703
rect 1176 -1288 1400 643
rect 2576 1540 2800 2603
rect 2576 1484 2660 1540
rect 2716 1484 2800 1540
rect 2576 -153 2800 1484
rect 2576 -209 2661 -153
rect 2717 -209 2800 -153
rect 2576 -1288 2800 -209
use CS_Switch_16x2  CS_Switch_16x2_0 ~/CS_DAC/Magic_gf180mcuD
timestamp 1755760707
transform 1 0 4010 0 1 -145
box -377 631 825 1384
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 74 0 1 725
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2874 0 -1 605
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  gf180mcu_fd_sc_mcu7t5v0__nand2_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 1514 0 -1 605
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 74 0 -1 605
box -86 -86 1206 870
<< labels >>
flabel metal1 206 149 278 402 1 FreeSans 800 0 0 0 Ri
port 1 n
flabel metal1 430 -73 502 319 1 FreeSans 800 0 0 0 Ci
port 2 n
flabel metal1 1638 181 2320 245 1 FreeSans 800 0 0 0 Ri-1
port 3 n
flabel metal1 204 1079 392 1155 1 FreeSans 800 0 0 0 CLK
port 4 n
flabel metal1 3973 1053 4029 1472 1 FreeSans 800 0 0 0 OUTP
port 5 n
rlabel metal1 3963 977 4039 1053 1 OUTP
port 5 n
flabel metal1 4455 1053 4511 1411 1 FreeSans 800 0 0 0 OUTN
port 6 n
rlabel metal1 4445 977 4521 1053 1 OUTN
port 6 n
flabel metal2 4423 -53 4479 837 1 FreeSans 800 0 0 0 VBIAS
port 7 n
rlabel metal2 4412 827 4488 903 1 VBIAS
port 7 n
flabel metal3 2576 -336 2800 1792 1 FreeSans 3200 0 0 0 VDD
port 8 n
flabel metal3 1176 -336 1400 1792 1 FreeSans 3200 0 0 0 VSS
port 9 n
rlabel metal3 1176 -1288 1400 -309 1 VSS
port 9 n
rlabel metal3 2576 -1288 2800 -309 1 VDD
port 8 n
rlabel metal3 1176 1624 1400 2603 1 VSS
port 9 n
rlabel metal3 2576 1624 2800 2603 1 VDD
port 8 n
<< end >>
