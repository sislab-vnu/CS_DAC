magic
tech gf180mcuD
magscale 1 10
timestamp 1758622075
<< nwell >>
rect 2999 1486 3100 1542
rect 1254 -265 2878 253
<< pwell >>
rect 4528 1077 5667 1239
rect 1170 253 3408 674
rect 4523 547 5667 1077
rect 4523 253 5730 547
<< psubdiff >>
rect 1275 698 1375 719
rect 1275 639 1295 698
rect 1359 639 1375 698
rect 1275 619 1375 639
rect 2844 694 2944 718
rect 2844 636 2859 694
rect 2930 636 2944 694
rect 2844 618 2944 636
<< nsubdiff >>
rect 84 1545 184 1559
rect 84 1479 102 1545
rect 171 1479 184 1545
rect 84 1459 184 1479
rect 2421 1536 2521 1559
rect 2421 1479 2447 1536
rect 2508 1479 2521 1536
rect 2421 1459 2521 1479
rect 1253 -151 1353 -131
rect 1253 -210 1274 -151
rect 1337 -210 1353 -151
rect 1253 -231 1353 -210
rect 2645 -160 2745 -127
rect 2645 -206 2673 -160
rect 2727 -206 2745 -160
rect 2645 -227 2745 -206
<< psubdiffcont >>
rect 1295 639 1359 698
rect 2859 636 2930 694
<< nsubdiffcont >>
rect 102 1479 171 1545
rect 2447 1479 2508 1536
rect 1274 -210 1337 -151
rect 2673 -206 2727 -160
<< metal1 >>
rect 204 1079 392 1155
rect 4868 1053 4924 1472
rect 5350 1053 5406 1411
rect 4858 977 4934 1053
rect 5340 977 5416 1053
rect 4891 893 5383 903
rect 4891 837 5318 893
rect 5374 837 5383 893
rect 4891 827 5383 837
rect 1191 639 1295 675
rect 1359 639 1530 675
rect 1191 545 1530 639
rect 2502 694 2928 714
rect 2502 636 2859 694
rect 2502 545 2928 636
rect 4426 545 4771 665
rect 206 149 278 402
rect 430 -73 502 319
rect 811 293 1638 350
rect 1638 181 2320 245
rect 1179 -151 1524 -119
rect 1179 -210 1274 -151
rect 1337 -210 1524 -151
rect 2514 -155 3198 -119
rect 1179 -239 1524 -210
rect 2514 -160 3010 -155
rect 2514 -206 2673 -160
rect 2727 -206 3010 -160
rect 2514 -211 3010 -206
rect 3111 -211 3198 -155
rect 2514 -239 3198 -211
<< via1 >>
rect 252 1478 364 1534
rect 1540 1486 1652 1542
rect 2999 1486 3100 1542
rect 4249 1130 4301 1182
rect 3291 1063 3343 1115
rect 3697 1063 3749 1115
rect 5033 1134 5089 1190
rect 5185 1134 5241 1190
rect 1000 985 1052 1037
rect 5318 837 5374 893
rect 896 615 1009 729
rect 2269 604 2380 716
rect 3719 616 3831 727
rect 1969 409 2021 461
rect 3141 196 3193 248
rect 3353 199 3405 251
rect 3695 199 3747 251
rect 4247 230 4299 282
rect 252 -201 364 -145
rect 1541 -214 1653 -158
rect 3010 -211 3111 -155
<< metal2 >>
rect 417 1854 4522 1986
rect 433 1638 4538 1770
rect 223 1534 392 1568
rect 223 1478 252 1534
rect 364 1478 392 1534
rect 223 1456 392 1478
rect 1472 1542 1726 1567
rect 1472 1486 1540 1542
rect 1652 1486 1726 1542
rect 1472 1456 1726 1486
rect 2937 1542 3161 1567
rect 2937 1486 2999 1542
rect 3100 1486 3161 1542
rect 2937 1456 3161 1486
rect 4240 1190 5099 1199
rect 4240 1182 5033 1190
rect 3112 1115 3776 1146
rect 4240 1130 4249 1182
rect 4301 1134 5033 1182
rect 5089 1134 5099 1190
rect 4301 1130 5099 1134
rect 4240 1119 5099 1130
rect 5175 1190 5251 1199
rect 5175 1134 5185 1190
rect 5241 1134 5251 1190
rect 975 1037 2064 1079
rect 975 985 1000 1037
rect 1052 985 2064 1037
rect 975 959 2064 985
rect 840 729 1079 754
rect 840 615 896 729
rect 1009 615 1079 729
rect 840 586 1079 615
rect 1944 500 2064 959
rect 3112 1063 3291 1115
rect 3343 1063 3697 1115
rect 3749 1063 3776 1115
rect 3112 1034 3776 1063
rect 2185 716 2465 767
rect 2185 604 2269 716
rect 2380 604 2465 716
rect 2185 560 2465 604
rect 1944 461 2088 500
rect 1944 409 1969 461
rect 2021 409 2088 461
rect 1944 392 2088 409
rect 3112 248 3262 1034
rect 3673 727 3902 763
rect 3673 616 3719 727
rect 3831 616 3902 727
rect 3673 575 3902 616
rect 5175 298 5251 1134
rect 4240 282 5251 298
rect 3112 196 3141 248
rect 3193 196 3262 248
rect 3112 181 3262 196
rect 3335 251 3760 280
rect 3335 199 3353 251
rect 3405 199 3695 251
rect 3747 199 3760 251
rect 4240 230 4247 282
rect 4299 230 5251 282
rect 4240 218 5251 230
rect 5307 893 5383 903
rect 5307 837 5318 893
rect 5374 837 5383 893
rect 3335 175 3760 199
rect 5307 -59 5383 837
rect 224 -145 393 -123
rect 224 -201 252 -145
rect 364 -201 393 -145
rect 224 -235 393 -201
rect 1487 -158 1712 -129
rect 1487 -214 1541 -158
rect 1653 -214 1712 -158
rect 1487 -233 1712 -214
rect 2968 -155 3168 -118
rect 2968 -211 3010 -155
rect 3111 -211 3168 -155
rect 2968 -224 3168 -211
<< via2 >>
rect 252 1478 364 1534
rect 1540 1486 1652 1542
rect 2999 1486 3100 1542
rect 896 615 1009 729
rect 2269 604 2380 716
rect 3719 616 3831 727
rect 252 -201 364 -145
rect 1541 -214 1653 -158
rect 3010 -211 3111 -155
<< metal3 >>
rect 140 1534 484 3283
rect 140 1478 252 1534
rect 364 1478 484 1534
rect 140 329 484 1478
rect 140 246 265 329
rect 357 246 484 329
rect 140 -145 484 246
rect 140 -201 252 -145
rect 364 -201 484 -145
rect 140 -852 484 -201
rect 789 929 1133 3283
rect 789 846 901 929
rect 993 846 1133 929
rect 789 729 1133 846
rect 789 615 896 729
rect 1009 615 1133 729
rect 789 -126 1133 615
rect 789 -218 890 -126
rect 1009 -218 1133 -126
rect 789 -850 1133 -218
rect 1432 1542 1776 3283
rect 1432 1486 1540 1542
rect 1652 1486 1776 1542
rect 1432 360 1776 1486
rect 1432 268 1533 360
rect 1652 268 1776 360
rect 1432 -158 1776 268
rect 1432 -214 1541 -158
rect 1653 -214 1776 -158
rect 1432 -857 1776 -214
rect 2159 936 2503 3277
rect 2159 853 2303 936
rect 2395 853 2503 936
rect 2159 716 2503 853
rect 2159 604 2269 716
rect 2380 604 2503 716
rect 2159 -120 2503 604
rect 2159 -212 2286 -120
rect 2405 -212 2503 -120
rect 2159 -850 2503 -212
rect 2889 1542 3233 3284
rect 2889 1486 2999 1542
rect 3100 1486 3233 1542
rect 2889 383 3233 1486
rect 2889 291 2987 383
rect 3106 291 3233 383
rect 2889 -155 3233 291
rect 2889 -211 3010 -155
rect 3111 -211 3233 -155
rect 2889 -856 3233 -211
rect 3614 981 3958 3269
rect 3614 898 3741 981
rect 3833 898 3958 981
rect 3614 727 3958 898
rect 3614 616 3719 727
rect 3831 616 3958 727
rect 3614 -129 3958 616
rect 3614 -221 3737 -129
rect 3856 -221 3958 -129
rect 3614 -850 3958 -221
<< via3 >>
rect 252 1478 364 1534
rect 265 246 357 329
rect 901 846 993 929
rect 890 -218 1009 -126
rect 1540 1486 1652 1542
rect 1533 268 1652 360
rect 2303 853 2395 936
rect 2286 -212 2405 -120
rect 2999 1486 3100 1542
rect 2987 291 3106 383
rect 3741 898 3833 981
rect 3737 -221 3856 -129
<< metal4 >>
rect -1095 1542 6313 1705
rect -1095 1534 1540 1542
rect -1095 1478 252 1534
rect 364 1486 1540 1534
rect 1652 1486 2999 1542
rect 3100 1486 6313 1542
rect 364 1478 6313 1486
rect -1095 1359 6313 1478
rect -1095 1358 -406 1359
rect -1114 981 6313 1065
rect -1114 936 3741 981
rect -1114 929 2303 936
rect -1114 846 901 929
rect 993 853 2303 929
rect 2395 898 3741 936
rect 3833 898 6313 981
rect 2395 853 6313 898
rect 993 846 6313 853
rect -1114 719 6313 846
rect -1114 718 -425 719
rect -1103 383 6332 478
rect -1103 360 2987 383
rect -1103 329 1533 360
rect -1103 246 265 329
rect 357 268 1533 329
rect 1652 291 2987 360
rect 3106 291 6332 383
rect 1652 268 6332 291
rect 357 246 6332 268
rect -1103 132 6332 246
rect -1103 131 -414 132
rect -1083 -63 -394 -62
rect -1083 -120 6338 -63
rect -1083 -126 2286 -120
rect -1083 -218 890 -126
rect 1009 -212 2286 -126
rect 2405 -129 6338 -120
rect 2405 -212 3737 -129
rect 1009 -218 3737 -212
rect -1083 -221 3737 -218
rect 3856 -221 6338 -129
rect -1083 -409 6338 -221
use CS_Switch_16x2  CS_Switch_16x2_0
timestamp 1755760707
transform 1 0 4905 0 1 -145
box -377 631 825 1384
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_1 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 3546 0 1 725
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_2
timestamp 1753044640
transform 1 0 3546 0 -1 605
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 74 0 1 725
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2874 0 -1 605
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  gf180mcu_fd_sc_mcu7t5v0__nand2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 1514 0 -1 605
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 74 0 -1 605
box -86 -86 1206 870
<< labels >>
flabel metal3 827 1749 1093 2241 1 FreeSans 800 0 0 0 VSS
port 9 n
flabel metal3 177 1774 443 2266 1 FreeSans 800 0 0 0 VDD
port 8 n
flabel metal1 204 1079 392 1155 1 FreeSans 400 0 0 0 CLK
port 4 n
flabel metal1 1638 181 2320 245 1 FreeSans 400 0 0 0 Ri-1
port 3 n
flabel metal1 430 -73 502 319 1 FreeSans 400 0 0 0 Ci
port 2 n
flabel metal1 206 149 278 402 1 FreeSans 400 0 0 0 Ri
port 1 n
flabel metal1 4872 1055 4922 1470 1 FreeSans 400 0 0 0 OUTP
port 5 n
flabel metal1 5353 1061 5402 1406 1 FreeSans 400 0 0 0 OUTN
port 6 n
flabel metal2 5321 -53 5371 820 1 FreeSans 400 0 0 0 VBIAS
port 7 n
<< end >>
