** sch_path: /home/ducluong/CS_DAC/xschem/test_symbols.sch
**.subckt test_symbols
x1 D3 CLK q1 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
x2 D2 CLK q2 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
x3 D CLK q4 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__dffq_4
V1 CLK GND PULSE(0 3.3 0 1n 1n 4n 10n)
V2 D GND PULSE(0 3.3 0 1n 1n 39n 80n)
V3 A1 GND PULSE(0 3.3 0 1n 1n 4n 10n)
V4 A2 GND PULSE(0 3.3 0 1n 1n 9n 20n)
x6 A1 A2 and1 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
x5 A1 A2 and4 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
x7 A1 i1 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x8 A1 i2 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
x9 A1 i3 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
x11 A1 A2 or1 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
x12 A1 A2 or2 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
x13 A1 A2 or4 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
x14 A1 A2 nand1 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
x15 A1 A2 nand2 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
x16 A1 A2 nand4 VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
V5 D2 GND PULSE(0 3.3 0 1n 1n 19n 40n)
V6 D3 GND PULSE(0 3.3 0 1n 1n 4n 10n)
x17 A1 A2 A3 nand3_1_zn VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__nand3_1
x18 A1 A2 A3 nor3_1_zn VDD VNW VPW VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
V7 A3 GND PULSE(0 3.3 0 1n 1n 50n 100n)
V8 VDD1 GND 3.3
x4 A1 A2 and2 VDD1 VDD1 GND GND gf180mcu_fd_sc_mcu7t5v0__or2_2
**** begin user architecture code

.include /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_typical
* .lib /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_statistical

 .include /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/spice/gf180mcu_fd_sc_mcu7t5v0.spice


.tran 1n 320n
.save all

**** end user architecture code
**.ends
.GLOBAL GND
.end
