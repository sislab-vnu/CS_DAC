magic
tech gf180mcuD
magscale 1 10
timestamp 1754903761
<< pwell >>
rect 426 1024 1804 1719
<< nmos >>
rect 496 1400 552 1444
rect 728 1400 784 1444
rect 956 1400 1012 1444
rect 1292 1366 1348 1478
rect 1440 1360 1500 1484
rect 1652 1360 1712 1484
<< ndiff >>
rect 602 1445 682 1462
rect 602 1444 619 1445
rect 450 1400 496 1444
rect 552 1400 619 1444
rect 602 1399 619 1400
rect 665 1444 682 1445
rect 830 1446 910 1462
rect 830 1444 846 1446
rect 665 1400 728 1444
rect 784 1400 846 1444
rect 665 1399 682 1400
rect 602 1382 682 1399
rect 830 1398 846 1400
rect 894 1444 910 1446
rect 1394 1478 1440 1484
rect 1246 1462 1292 1478
rect 1058 1445 1138 1462
rect 1058 1444 1075 1445
rect 894 1400 956 1444
rect 1012 1400 1075 1444
rect 894 1398 910 1400
rect 830 1382 910 1398
rect 1058 1399 1075 1400
rect 1121 1399 1138 1445
rect 1058 1382 1138 1399
rect 1198 1446 1292 1462
rect 1198 1398 1214 1446
rect 1262 1398 1292 1446
rect 1198 1382 1292 1398
rect 1246 1366 1292 1382
rect 1348 1366 1440 1478
rect 1394 1360 1440 1366
rect 1500 1462 1546 1484
rect 1606 1462 1652 1484
rect 1500 1446 1652 1462
rect 1500 1398 1532 1446
rect 1580 1398 1652 1446
rect 1500 1382 1652 1398
rect 1500 1360 1546 1382
rect 1606 1360 1652 1382
rect 1712 1360 1758 1484
<< ndiffc >>
rect 619 1399 665 1445
rect 846 1398 894 1446
rect 1075 1399 1121 1445
rect 1214 1398 1262 1446
rect 1532 1398 1580 1446
<< polysilicon >>
rect 716 1553 796 1570
rect 716 1507 733 1553
rect 779 1507 796 1553
rect 716 1490 796 1507
rect 944 1553 1024 1570
rect 944 1507 961 1553
rect 1007 1507 1024 1553
rect 944 1490 1024 1507
rect 1292 1568 1500 1581
rect 1292 1522 1350 1568
rect 1450 1522 1500 1568
rect 1292 1504 1500 1522
rect 496 1444 552 1490
rect 496 1354 552 1400
rect 728 1444 784 1490
rect 728 1354 784 1400
rect 956 1444 1012 1490
rect 1292 1478 1348 1504
rect 1440 1484 1500 1504
rect 1652 1484 1712 1528
rect 956 1354 1012 1400
rect 488 1341 560 1354
rect 488 1295 501 1341
rect 547 1295 560 1341
rect 1292 1320 1348 1366
rect 1440 1314 1500 1360
rect 1652 1314 1712 1360
rect 488 1282 560 1295
rect 1646 1301 1718 1314
rect 1646 1255 1659 1301
rect 1705 1255 1718 1301
rect 1646 1242 1718 1255
<< polycontact >>
rect 733 1507 779 1553
rect 961 1507 1007 1553
rect 1350 1522 1450 1568
rect 501 1295 547 1341
rect 1659 1255 1705 1301
<< metal1 >>
rect 1315 1568 1478 1576
rect 718 1553 794 1568
rect 718 1507 733 1553
rect 779 1507 794 1553
rect 718 1492 794 1507
rect 946 1553 1022 1568
rect 946 1507 961 1553
rect 1007 1507 1022 1553
rect 1315 1522 1350 1568
rect 1450 1522 1478 1568
rect 1315 1512 1478 1522
rect 946 1492 1022 1507
rect 604 1445 680 1460
rect 604 1399 619 1445
rect 665 1399 680 1445
rect 604 1384 680 1399
rect 832 1446 908 1460
rect 832 1398 846 1446
rect 894 1398 908 1446
rect 832 1384 908 1398
rect 1060 1445 1136 1460
rect 1060 1399 1075 1445
rect 1121 1399 1136 1445
rect 1060 1384 1136 1399
rect 1200 1446 1276 1460
rect 1200 1398 1214 1446
rect 1262 1398 1276 1446
rect 1200 1384 1276 1398
rect 1518 1446 1594 1460
rect 1518 1398 1532 1446
rect 1580 1398 1594 1446
rect 1518 1384 1594 1398
rect 501 1341 547 1352
rect 501 1231 547 1295
rect 846 1332 894 1384
rect 1214 1332 1262 1384
rect 846 1284 1262 1332
rect 1152 1283 1262 1284
rect 1532 1231 1580 1384
rect 1659 1301 1705 1312
rect 1659 1231 1705 1255
rect 458 1120 1796 1231
<< labels >>
flabel metal1 1315 1512 1478 1576 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel pwell 619 1123 734 1226 1 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
flabel metal1 784 1120 1624 1231 1 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional
flabel metal1 718 1492 794 1568 1 FreeSans 400 0 0 0 INP
port 1 n
flabel metal1 946 1492 1022 1568 1 FreeSans 400 0 0 0 INN
port 2 n
flabel metal1 604 1384 680 1460 1 FreeSans 400 0 0 0 OUTP
port 3 n
flabel metal1 1060 1384 1136 1460 1 FreeSans 400 0 0 0 OUTN
port 4 n
<< end >>
