magic
tech gf180mcuD
magscale 1 10
timestamp 1755930310
<< metal1 >>
rect 11162 40089 11982 40395
rect 11162 39838 11423 40089
rect 11744 39838 11982 40089
rect 11162 39568 11982 39838
rect 11427 38589 11763 39568
rect 38229 39387 39060 39637
rect 38229 39076 38473 39387
rect 38774 39076 39060 39387
rect 38229 38817 39060 39076
rect 11426 35831 11764 38589
rect 38373 37641 38913 38817
rect 11423 35744 11764 35831
rect 11423 32986 11761 35744
rect 38374 33096 38912 37641
rect 38370 33022 38912 33096
rect 11424 26544 11760 32986
rect 38370 28639 38910 33022
rect 33884 28567 38910 28639
rect 33882 28099 38910 28567
rect 33882 27642 34176 28099
rect 47920 28056 54417 28058
rect 41274 28052 54417 28056
rect 41274 27532 54430 28052
rect 41274 27530 48003 27532
rect 25536 26742 25872 26880
rect 25536 26686 25676 26742
rect 25732 26686 25872 26742
rect 25536 26544 25872 26686
rect 11480 25928 11704 26544
rect -952 25592 11704 25928
rect -952 20425 -615 25592
rect 9799 25370 10404 25371
rect 13247 25370 14416 25372
rect 25592 25370 25816 26544
rect 53901 26369 54430 27532
rect 53438 25894 54902 26369
rect 53438 25401 53838 25894
rect 54471 25401 54902 25894
rect -392 25034 29848 25370
rect -392 25033 11497 25034
rect 12181 25033 29848 25034
rect -316 24043 -221 25033
rect -133 24829 -37 24925
rect -133 24774 -112 24829
rect -56 24774 -37 24829
rect -133 24293 -37 24774
rect -317 23882 -221 24043
rect -132 24041 -37 24293
rect 8287 24152 8395 25033
rect 8287 24085 8300 24152
rect 8381 24085 8395 24152
rect 8287 24071 8395 24085
rect 18009 24128 18091 25033
rect 18009 24076 18021 24128
rect 18079 24076 18091 24128
rect 28146 24178 28216 25033
rect 53438 24945 54902 25401
rect 28146 24122 28151 24178
rect 28207 24122 28216 24178
rect 28146 24108 28216 24122
rect -133 23969 -37 24041
rect -317 23614 -222 23882
rect -133 23788 -38 23969
rect -133 23707 -37 23788
rect 33880 23761 34159 24481
rect -318 23420 -222 23614
rect -318 23147 -223 23420
rect -132 23261 -37 23707
rect 28147 23572 28213 23586
rect 18014 23527 18085 23539
rect -132 23166 309 23261
rect 8287 23236 8395 23300
rect -132 23165 -37 23166
rect -318 22991 -221 23147
rect 8287 23168 8307 23236
rect 8379 23168 8395 23236
rect -316 22753 -221 22991
rect -317 22524 -221 22753
rect 8287 22819 8395 23168
rect 8589 23243 9036 23274
rect 8589 23169 8680 23243
rect 8793 23169 9036 23243
rect 8589 23154 9036 23169
rect 13825 23240 15130 23274
rect 13825 23184 13888 23240
rect 13944 23184 15130 23240
rect 13825 23154 15130 23184
rect 8287 22721 9191 22819
rect 18014 22800 18085 23471
rect 28147 23520 28155 23572
rect 28208 23520 28213 23572
rect 18192 23240 18753 23274
rect 18192 23184 18283 23240
rect 18339 23184 18753 23240
rect 18192 23154 18753 23184
rect 23438 23240 24803 23274
rect 23438 23184 23493 23240
rect 23549 23184 24803 23240
rect 23438 23154 24803 23184
rect 28147 22852 28213 23520
rect 29296 23154 29448 23274
rect 18014 22729 18820 22800
rect 28147 22786 28508 22852
rect 41270 22768 41608 24364
rect 8287 22720 8395 22721
rect -317 22225 -222 22524
rect 11045 22465 11946 22491
rect 11045 22389 11761 22465
rect 11874 22389 11946 22465
rect 11045 22369 11946 22389
rect 15764 22456 16758 22490
rect 15764 22400 16605 22456
rect 16661 22400 16758 22456
rect 15764 22368 16758 22400
rect 20732 22456 21585 22490
rect 20732 22400 21421 22456
rect 21477 22400 21585 22456
rect 20732 22370 21585 22400
rect 25777 22456 26400 22490
rect 25777 22400 26292 22456
rect 26348 22400 26400 22456
rect 25777 22370 26400 22400
rect 30382 22456 31263 22490
rect 30382 22400 31111 22456
rect 31167 22400 31263 22456
rect 30382 22370 31263 22400
rect -317 22130 306 22225
rect -952 20350 307 20425
rect -952 15780 -615 20350
rect 6040 19995 6311 20115
rect 6042 17195 6313 17315
rect -952 15721 287 15780
rect -952 10248 -615 15721
rect 5995 14395 6266 14515
rect 6832 13374 7056 13403
rect 6832 13305 6885 13374
rect 7001 13305 7056 13374
rect 6832 13283 7056 13305
rect 6046 11595 6317 11715
rect -952 10180 297 10248
rect -952 4582 -615 10180
rect 27833 9733 28055 9762
rect 27833 9663 27888 9733
rect 28000 9663 28055 9733
rect 27833 9634 28055 9663
rect 6046 8795 6317 8915
rect 27831 6939 28053 6967
rect 27831 6869 27887 6939
rect 27999 6869 28053 6939
rect 27831 6832 28053 6869
rect 6047 5995 6318 6115
rect -952 4521 330 4582
rect -952 2800 -615 4521
rect 6052 3195 6323 3315
rect 6043 395 6314 515
<< via1 >>
rect 11423 39838 11744 40089
rect 38473 39076 38774 39387
rect 35784 27796 35874 27869
rect 37124 27023 37213 27079
rect 35801 26846 35890 26918
rect 25676 26686 25732 26742
rect 37123 26063 37244 26128
rect 35794 25881 35883 25953
rect 53838 25401 54471 25894
rect 37126 25104 37244 25163
rect -112 24774 -56 24829
rect 8300 24085 8381 24152
rect 18021 24076 18079 24128
rect 35800 24915 35893 24993
rect 28151 24122 28207 24178
rect 37119 24130 37237 24189
rect 18014 23471 18085 23527
rect 470 23133 526 23187
rect 8307 23168 8379 23236
rect 8680 23169 8793 23243
rect 13888 23184 13944 23240
rect 391 22657 504 22733
rect 9350 22790 9409 22850
rect 10361 22794 10415 22848
rect 15127 22763 15182 22816
rect 28155 23520 28208 23572
rect 18283 23184 18339 23240
rect 23493 23184 23549 23240
rect 28442 23177 28542 23245
rect 18982 22794 19043 22850
rect 20104 22792 20160 22848
rect 24918 22793 24979 22852
rect 25144 22792 25200 22848
rect 28671 22793 28732 22850
rect 29788 22792 29852 22852
rect 3881 22614 3971 22672
rect 11761 22389 11874 22465
rect 16605 22400 16661 22456
rect 21421 22400 21477 22456
rect 26292 22400 26348 22456
rect 31111 22400 31167 22456
rect 4090 22229 4144 22282
rect 3865 22172 3920 22224
rect 2184 21703 2296 21777
rect 6887 21698 7001 21776
rect 11760 21700 11873 21782
rect 16593 21710 16683 21769
rect 21412 21709 21490 21773
rect 26264 21706 26375 21776
rect 31080 21714 31193 21771
rect 37146 21707 37224 21773
rect 244 21380 302 21434
rect 470 21325 525 21377
rect 392 20849 505 20925
rect 3864 20871 3976 20940
rect 8678 20855 8793 20940
rect 13889 20866 14003 20934
rect 18268 20864 18348 20943
rect 23462 20862 23576 20944
rect 27887 20864 28000 20937
rect 33039 20874 33155 20938
rect 35784 20869 35896 20928
rect 2184 20019 2296 20085
rect 6888 20014 7000 20091
rect 11760 20016 11872 20098
rect 16583 20022 16673 20081
rect 21409 20021 21486 20085
rect 26277 20017 26366 20089
rect 31079 20020 31192 20077
rect 37145 20023 37223 20089
rect 2184 18907 2296 18973
rect 6888 18901 7000 18976
rect 11760 18904 11872 18986
rect 16593 18910 16665 18969
rect 21404 18914 21481 18978
rect 26281 18903 26370 18975
rect 31080 18911 31192 18969
rect 37151 18909 37227 18978
rect 392 18005 505 18072
rect 3863 18059 3977 18136
rect 8680 18055 8792 18139
rect 13888 18070 14002 18138
rect 18269 18065 18349 18144
rect 23464 18068 23575 18143
rect 27889 18066 28002 18139
rect 33038 18053 33154 18117
rect 35784 18068 35896 18127
rect 454 17621 510 17673
rect 231 17561 284 17616
rect 2184 17214 2296 17300
rect 6888 17221 7000 17291
rect 11761 17212 11872 17282
rect 16599 17219 16671 17278
rect 21407 17212 21487 17285
rect 26270 17214 26369 17285
rect 31080 17221 31192 17279
rect 37143 17220 37219 17289
rect 2184 16117 2296 16181
rect 6887 16104 7000 16173
rect 11762 16110 11873 16180
rect 16588 16114 16667 16175
rect 21411 16108 21491 16181
rect 26271 16105 26370 16176
rect 31080 16115 31192 16171
rect 37144 16111 37218 16175
rect 450 15724 505 15779
rect 378 15254 513 15321
rect 3863 15255 3977 15332
rect 8679 15249 8791 15343
rect 13887 15263 14008 15338
rect 18267 15261 18351 15336
rect 23462 15258 23577 15324
rect 27888 15263 28000 15334
rect 33040 15269 33152 15339
rect 35784 15274 35896 15333
rect 224 14765 280 14819
rect 2184 14425 2296 14495
rect 6888 14420 7001 14489
rect 11760 14418 11873 14494
rect 16592 14417 16671 14478
rect 21397 14410 21484 14481
rect 26265 14414 26371 14483
rect 31080 14423 31192 14479
rect 37150 14425 37224 14489
rect 2184 13310 2296 13383
rect 6885 13305 7001 13374
rect 11760 13308 11873 13384
rect 16594 13308 16668 13372
rect 21406 13305 21493 13376
rect 26267 13311 26373 13380
rect 31080 13310 31192 13370
rect 37148 13308 37226 13376
rect 3864 12464 3977 12535
rect 396 12402 501 12463
rect 8681 12455 8793 12549
rect 13885 12460 14006 12535
rect 18268 12455 18352 12530
rect 23462 12460 23577 12526
rect 27889 12456 28001 12527
rect 33040 12465 33152 12535
rect 35784 12465 35896 12524
rect 450 11987 507 12043
rect 2184 11616 2296 11700
rect 6886 11615 7002 11684
rect 11760 11611 11872 11686
rect 16601 11617 16675 11681
rect 21397 11610 21483 11686
rect 26278 11611 26367 11687
rect 31080 11625 31192 11685
rect 37146 11618 37224 11686
rect 2184 10503 2296 10581
rect 6887 10505 7001 10576
rect 11760 10508 11872 10583
rect 16593 10512 16669 10574
rect 21402 10500 21488 10576
rect 26277 10506 26366 10582
rect 31080 10518 31193 10573
rect 37137 10506 37219 10579
rect 461 10123 516 10178
rect 368 9654 474 9719
rect 3863 9670 3976 9741
rect 8680 9647 8794 9730
rect 13887 9663 14004 9735
rect 18265 9655 18353 9735
rect 23463 9663 23578 9726
rect 27888 9663 28000 9733
rect 33031 9666 33143 9732
rect 35784 9674 35896 9732
rect 347 9217 404 9274
rect 2184 8813 2296 8893
rect 6886 8814 7000 8885
rect 11760 8811 11872 8889
rect 16598 8816 16674 8878
rect 21397 8811 21484 8885
rect 26265 8811 26364 8886
rect 31079 8826 31192 8882
rect 37142 8812 37224 8885
rect 2184 7714 2296 7784
rect 6888 7708 7000 7773
rect 11760 7703 11872 7781
rect 16589 7706 16670 7772
rect 21404 7705 21491 7779
rect 26273 7708 26372 7783
rect 31079 7716 31192 7772
rect 37144 7711 37228 7779
rect 390 6805 505 6874
rect 3863 6854 3977 6935
rect 8679 6849 8791 6928
rect 13886 6866 14003 6938
rect 18263 6876 18351 6956
rect 23462 6865 23577 6928
rect 27887 6869 27999 6939
rect 33041 6864 33153 6930
rect 35784 6863 35896 6921
rect 334 6421 389 6473
rect 554 6416 618 6479
rect 2184 6012 2296 6088
rect 6888 6016 7000 6081
rect 11761 6016 11874 6089
rect 16593 6016 16674 6082
rect 21400 6011 21485 6083
rect 26275 6010 26367 6090
rect 31080 6026 31193 6082
rect 37140 6015 37224 6083
rect 2184 4910 2296 4984
rect 6888 4903 7001 4974
rect 11759 4907 11872 4980
rect 16589 4906 16672 4976
rect 21408 4902 21493 4974
rect 26281 4900 26373 4980
rect 31080 4921 31192 4977
rect 37140 4910 37228 4976
rect 557 4523 611 4577
rect 390 4062 507 4141
rect 3863 4058 3977 4139
rect 8680 4052 8793 4129
rect 13887 4060 14000 4135
rect 18267 4066 18360 4141
rect 23460 4056 23576 4127
rect 27887 4050 28001 4123
rect 33030 4072 33139 4136
rect 35783 4074 35896 4130
rect 333 3620 388 3674
rect 2184 3214 2296 3293
rect 6888 3217 7001 3288
rect 11757 3209 11875 3284
rect 16594 3218 16677 3288
rect 21401 3212 21486 3283
rect 26264 3210 26360 3290
rect 31080 3222 31192 3278
rect 37137 3219 37225 3285
rect 2184 2104 2296 2172
rect 6887 2104 7001 2173
rect 11758 2106 11876 2181
rect 16595 2104 16675 2177
rect 21403 2103 21488 2174
rect 26276 2099 26372 2179
rect 31079 2117 31193 2178
rect 3864 1265 3976 1332
rect 8679 1257 8792 1334
rect 13872 1255 14002 1328
rect 18262 1260 18355 1335
rect 23462 1271 23578 1342
rect 27887 1257 28001 1330
rect 33043 1265 33152 1329
rect 2184 416 2296 489
rect 6887 418 7001 487
rect 11760 410 11872 487
rect 16588 412 16668 485
rect 21402 408 21481 480
rect 26275 406 26363 483
rect 31079 421 31193 482
<< metal2 >>
rect 3166 39659 3986 40486
rect 3419 38742 3757 39659
rect 8115 39645 8935 40472
rect 11162 40089 11982 40395
rect 11162 39838 11423 40089
rect 11744 39838 11982 40089
rect 3416 37641 3757 38742
rect 8347 38561 8683 39645
rect 11162 39568 11982 39838
rect 16947 39645 17767 40472
rect 21605 39810 22425 40637
rect 25302 39863 26122 40690
rect 31082 40348 31902 41179
rect 8339 37641 8683 38561
rect 17194 38076 17530 39645
rect 17194 37641 17534 38076
rect 21843 38057 22179 39810
rect 3416 33276 3754 37641
rect 8339 35838 8677 37641
rect 8339 35716 8680 35838
rect 3414 26767 3758 33276
rect 8342 32993 8680 35716
rect 17196 35369 17534 37641
rect 3414 26656 3528 26767
rect 3640 26656 3758 26767
rect 3414 26543 3758 26656
rect 8344 26544 8680 32993
rect 17190 35231 17534 35369
rect 21841 37641 22179 38057
rect 25539 37998 25875 39863
rect 31232 38941 31568 40348
rect 32703 39616 33523 40447
rect 34952 39980 35772 40811
rect 36320 39983 37140 40814
rect 31229 38062 31568 38941
rect 25539 37641 25877 37998
rect 17190 26707 17528 35231
rect 21841 33096 22169 37641
rect 25549 33096 25877 37641
rect 31228 37641 31568 38062
rect 32927 37641 33263 39616
rect 35163 38027 35499 39980
rect 35152 37641 35499 38027
rect 36545 37957 36881 39983
rect 38229 39387 39060 39637
rect 38229 39076 38473 39387
rect 38774 39076 39060 39387
rect 38229 38817 39060 39076
rect 36545 37656 36885 37957
rect 36549 37641 36885 37656
rect 31228 33096 31556 37641
rect 32930 33096 33258 37641
rect 35152 33096 35480 37641
rect 36550 33096 36878 37641
rect 17190 26600 17300 26707
rect 17418 26600 17528 26707
rect 17190 26544 17528 26600
rect 21840 26544 22176 33096
rect 25536 32940 25877 33096
rect 25536 26742 25872 32940
rect 25536 26686 25676 26742
rect 25732 26686 25872 26742
rect 25536 26544 25872 26686
rect 31226 27429 31565 33096
rect 8400 26376 8625 26544
rect -1344 26371 8625 26376
rect -1344 26040 8624 26371
rect -1344 21444 -1007 26040
rect 11535 24977 12172 24978
rect 21896 24977 22120 26544
rect 31226 25709 31562 27429
rect 32924 26661 33260 33096
rect 35152 32969 35496 33096
rect 35160 27297 35496 32969
rect 35755 27869 35905 27885
rect 35755 27796 35784 27869
rect 35874 27796 35905 27869
rect 35755 27786 35905 27796
rect 35768 26918 35918 26931
rect 35768 26846 35801 26918
rect 35890 26846 35918 26918
rect 35768 26832 35918 26846
rect 32924 26555 35399 26661
rect 32928 26327 35399 26555
rect 35772 25953 35906 25968
rect 35772 25881 35794 25953
rect 35883 25881 35906 25953
rect 35772 25873 35906 25881
rect 31226 25369 35417 25709
rect 35790 24993 35903 25003
rect -168 24829 30070 24977
rect 35790 24915 35800 24993
rect 35893 24915 35903 24993
rect 35790 24905 35903 24915
rect -168 24774 -112 24829
rect -56 24774 30070 24829
rect -168 24641 30070 24774
rect 36546 24719 36882 33096
rect 52171 30107 53635 31531
rect 40270 29352 46999 29353
rect 52638 29352 53162 30107
rect 40270 29131 53162 29352
rect 40270 29049 40384 29131
rect 40502 29049 53162 29131
rect 40270 28831 53162 29049
rect 40270 28827 53157 28831
rect 46660 28826 53157 28827
rect 55903 28710 57367 29206
rect 40770 28707 47499 28709
rect 53727 28707 57367 28710
rect 40770 28183 57367 28707
rect 40770 28048 41101 28183
rect 47315 28181 57367 28183
rect 53727 28179 57367 28181
rect 55903 27782 57367 28179
rect 37091 27079 37246 27100
rect 37091 27023 37124 27079
rect 37213 27023 37246 27079
rect 37091 27004 37246 27023
rect 37106 26128 37262 26143
rect 37106 26063 37123 26128
rect 37244 26063 37262 26128
rect 37106 26050 37262 26063
rect 53438 25894 54902 26369
rect 53438 25401 53838 25894
rect 54471 25401 54902 25894
rect 37106 25163 37262 25179
rect 37106 25104 37126 25163
rect 37244 25104 37262 25163
rect 37106 25086 37262 25104
rect 53438 24945 54902 25401
rect -168 24640 13276 24641
rect 14319 24640 30070 24641
rect 453 24380 548 24499
rect 453 24324 472 24380
rect 530 24324 548 24380
rect 453 23187 548 24324
rect 453 23133 470 23187
rect 526 23133 548 23187
rect 453 23121 548 23133
rect 336 22733 562 22762
rect 336 22657 391 22733
rect 504 22657 562 22733
rect 336 22628 562 22657
rect 3836 22672 4021 22707
rect 3836 22614 3881 22672
rect 3971 22614 4021 22672
rect 3836 22586 4021 22614
rect 4080 22292 4152 24640
rect 8287 24152 8395 24160
rect 8287 24085 8300 24152
rect 8381 24085 8395 24152
rect 8287 23258 8395 24085
rect 8272 23236 8403 23258
rect 8272 23168 8307 23236
rect 8379 23168 8403 23236
rect 8272 23148 8403 23168
rect 8624 23243 8847 23275
rect 8624 23169 8680 23243
rect 8793 23169 8847 23243
rect 8624 23154 8847 23169
rect 9342 22857 9414 24640
rect 13878 23240 13954 23250
rect 13878 23184 13888 23240
rect 13944 23184 13954 23240
rect 13878 23174 13954 23184
rect 9327 22850 9428 22857
rect 9327 22790 9350 22850
rect 9409 22790 9428 22850
rect 9327 22785 9428 22790
rect 10348 22850 10428 22860
rect 10348 22792 10358 22850
rect 10418 22792 10428 22850
rect 15121 22828 15185 24640
rect 18014 24128 18085 24140
rect 18014 24076 18021 24128
rect 18079 24076 18085 24128
rect 18014 23541 18085 24076
rect 17999 23527 18095 23541
rect 17999 23471 18014 23527
rect 18085 23471 18095 23527
rect 17999 23462 18095 23471
rect 18273 23240 18349 23250
rect 18273 23184 18283 23240
rect 18339 23184 18349 23240
rect 18273 23174 18349 23184
rect 18976 22856 19048 24640
rect 20094 24416 20166 24426
rect 20094 24360 20104 24416
rect 20160 24360 20166 24416
rect 18968 22850 19057 22856
rect 10348 22782 10428 22792
rect 15114 22816 15195 22828
rect 15114 22763 15127 22816
rect 15182 22763 15195 22816
rect 18968 22794 18982 22850
rect 19043 22794 19057 22850
rect 18968 22788 19057 22794
rect 20094 22848 20166 24360
rect 23483 23240 23559 23250
rect 23483 23184 23493 23240
rect 23549 23184 23559 23240
rect 23483 23174 23559 23184
rect 24912 22860 24984 24640
rect 25134 24416 25206 24425
rect 25134 24360 25144 24416
rect 25200 24360 25206 24416
rect 20094 22792 20104 22848
rect 20160 22792 20166 22848
rect 20094 22780 20166 22792
rect 24905 22852 24993 22860
rect 24905 22793 24918 22852
rect 24979 22793 24993 22852
rect 24905 22785 24993 22793
rect 25134 22848 25206 24360
rect 28137 24178 28222 24185
rect 28137 24124 28151 24178
rect 28147 24122 28151 24124
rect 28207 24124 28222 24178
rect 28207 24122 28213 24124
rect 28147 23582 28213 24122
rect 28133 23572 28228 23582
rect 28133 23520 28155 23572
rect 28208 23520 28228 23572
rect 28133 23509 28228 23520
rect 27833 23261 28448 23262
rect 27833 23260 28553 23261
rect 27833 23251 28555 23260
rect 27833 23179 27862 23251
rect 28000 23245 28555 23251
rect 28000 23179 28442 23245
rect 27833 23177 28442 23179
rect 28542 23177 28555 23245
rect 27833 23167 28555 23177
rect 27938 23166 28555 23167
rect 28427 23164 28555 23166
rect 28662 22855 28734 24640
rect 35172 24382 36885 24719
rect 37086 24189 37271 24207
rect 37086 24130 37119 24189
rect 37237 24130 37271 24189
rect 37086 24118 37271 24130
rect 25134 22792 25144 22848
rect 25200 22792 25206 22848
rect 25134 22780 25206 22792
rect 28648 22850 28750 22855
rect 28648 22793 28671 22850
rect 28732 22793 28750 22850
rect 28648 22784 28750 22793
rect 29778 22852 29862 22862
rect 29778 22792 29788 22852
rect 29852 22792 29862 22852
rect 29778 22782 29862 22792
rect 40765 22781 41103 24377
rect 15114 22752 15195 22763
rect 11727 22465 11904 22491
rect 11727 22389 11761 22465
rect 11874 22389 11904 22465
rect 16595 22456 16671 22466
rect 16595 22400 16605 22456
rect 16661 22400 16671 22456
rect 16595 22390 16671 22400
rect 21411 22456 21487 22466
rect 21411 22400 21421 22456
rect 21477 22400 21487 22456
rect 21411 22390 21487 22400
rect 26282 22456 26358 22466
rect 26282 22400 26292 22456
rect 26348 22400 26358 22456
rect 26282 22390 26358 22400
rect 31101 22456 31177 22466
rect 31101 22400 31111 22456
rect 31167 22400 31177 22456
rect 31101 22390 31177 22400
rect 11727 22369 11904 22389
rect 4067 22282 4162 22292
rect 3851 22226 3934 22237
rect 3851 22170 3862 22226
rect 3923 22170 3934 22226
rect 4067 22229 4090 22282
rect 4144 22229 4162 22282
rect 4067 22213 4162 22229
rect 3851 22159 3934 22170
rect 2128 21777 2352 21803
rect 2128 21703 2184 21777
rect 2296 21703 2352 21777
rect 2128 21683 2352 21703
rect 6832 21776 7056 21803
rect 6832 21698 6887 21776
rect 7001 21698 7056 21776
rect 6832 21683 7056 21698
rect 11704 21782 11928 21803
rect 11704 21700 11760 21782
rect 11873 21700 11928 21782
rect 11704 21683 11928 21700
rect 16520 21769 16744 21803
rect 16520 21710 16593 21769
rect 16683 21710 16744 21769
rect 16520 21683 16744 21710
rect 21358 21773 21543 21792
rect 21358 21709 21412 21773
rect 21490 21709 21543 21773
rect 21358 21696 21543 21709
rect 26222 21776 26412 21792
rect 26222 21706 26264 21776
rect 26375 21706 26412 21776
rect 26222 21687 26412 21706
rect 31024 21771 31248 21792
rect 31024 21714 31080 21771
rect 31193 21714 31248 21771
rect 31024 21691 31248 21714
rect 37107 21773 37270 21793
rect 37107 21707 37146 21773
rect 37224 21707 37270 21773
rect 37107 21692 37270 21707
rect 230 21444 320 21449
rect -1344 21434 320 21444
rect -1344 21380 244 21434
rect 302 21380 320 21434
rect -1344 21376 320 21380
rect -1344 17545 -1007 21376
rect 230 21372 320 21376
rect 457 21380 538 21390
rect 457 21323 467 21380
rect 528 21323 538 21380
rect 457 21313 538 21323
rect 335 20925 559 20947
rect 335 20849 392 20925
rect 505 20849 559 20925
rect 335 20829 559 20849
rect 3808 20940 4034 20970
rect 3808 20871 3864 20940
rect 3976 20871 4034 20940
rect 3808 20844 4034 20871
rect 8623 20940 8848 20987
rect 8623 20855 8678 20940
rect 8793 20855 8848 20940
rect 8623 20822 8848 20855
rect 13856 20934 14035 20958
rect 13856 20866 13889 20934
rect 14003 20866 14035 20934
rect 13856 20835 14035 20866
rect 18231 20943 18383 20974
rect 18231 20864 18268 20943
rect 18348 20864 18383 20943
rect 18231 20834 18383 20864
rect 23408 20944 23632 20973
rect 23408 20862 23462 20944
rect 23576 20862 23632 20944
rect 23408 20832 23632 20862
rect 27831 20937 28057 20949
rect 27831 20864 27887 20937
rect 28000 20864 28057 20937
rect 27831 20833 28057 20864
rect 32984 20938 33208 20974
rect 32984 20874 33039 20938
rect 33155 20874 33208 20938
rect 32984 20848 33208 20874
rect 35736 20928 35937 20948
rect 35736 20869 35784 20928
rect 35896 20869 35937 20928
rect 35736 20845 35937 20869
rect 2128 20085 2352 20115
rect 2128 20019 2184 20085
rect 2296 20019 2352 20085
rect 2128 19995 2352 20019
rect 6832 20091 7057 20115
rect 6832 20014 6888 20091
rect 7000 20014 7057 20091
rect 6832 19995 7057 20014
rect 11704 20098 11928 20115
rect 11704 20016 11760 20098
rect 11872 20016 11928 20098
rect 11704 19995 11928 20016
rect 16540 20081 16720 20096
rect 16540 20022 16583 20081
rect 16673 20022 16720 20081
rect 16540 20004 16720 20022
rect 21355 20085 21540 20098
rect 21355 20021 21409 20085
rect 21486 20021 21540 20085
rect 21355 20006 21540 20021
rect 26228 20089 26418 20104
rect 26228 20017 26277 20089
rect 26366 20017 26418 20089
rect 26228 19999 26418 20017
rect 31023 20077 31248 20097
rect 31023 20020 31079 20077
rect 31192 20020 31248 20077
rect 31023 20003 31248 20020
rect 37092 20089 37277 20108
rect 37092 20023 37145 20089
rect 37223 20023 37277 20089
rect 37092 20006 37277 20023
rect 2128 18973 2352 19003
rect 2128 18907 2184 18973
rect 2296 18907 2352 18973
rect 2128 18883 2352 18907
rect 6832 18976 7056 19002
rect 6832 18901 6888 18976
rect 7000 18901 7056 18976
rect 6832 18883 7056 18901
rect 11704 18986 11928 19002
rect 11704 18904 11760 18986
rect 11872 18904 11928 18986
rect 11704 18883 11928 18904
rect 16540 18969 16720 18988
rect 16540 18910 16593 18969
rect 16665 18910 16720 18969
rect 16540 18896 16720 18910
rect 21371 18978 21516 18995
rect 21371 18914 21404 18978
rect 21481 18914 21516 18978
rect 21371 18897 21516 18914
rect 26221 18975 26417 18991
rect 26221 18903 26281 18975
rect 26370 18903 26417 18975
rect 26221 18887 26417 18903
rect 31024 18969 31249 18988
rect 31024 18911 31080 18969
rect 31192 18911 31249 18969
rect 31024 18894 31249 18911
rect 37099 18978 37284 18996
rect 37099 18909 37151 18978
rect 37227 18909 37284 18978
rect 37099 18894 37284 18909
rect 3807 18136 4033 18157
rect 336 18072 560 18097
rect 336 18005 392 18072
rect 505 18005 560 18072
rect 3807 18059 3863 18136
rect 3977 18059 4033 18136
rect 3807 18031 4033 18059
rect 8625 18139 8848 18176
rect 8625 18055 8680 18139
rect 8792 18055 8848 18139
rect 8625 18028 8848 18055
rect 13840 18138 14050 18175
rect 13840 18070 13888 18138
rect 14002 18070 14050 18138
rect 13840 18039 14050 18070
rect 18228 18144 18387 18174
rect 18228 18065 18269 18144
rect 18349 18065 18387 18144
rect 18228 18041 18387 18065
rect 23408 18143 23632 18167
rect 23408 18068 23464 18143
rect 23575 18068 23632 18143
rect 23408 18032 23632 18068
rect 27833 18139 28057 18167
rect 27833 18066 27889 18139
rect 28002 18066 28057 18139
rect 27833 18031 28057 18066
rect 32985 18117 33201 18139
rect 32985 18053 33038 18117
rect 33154 18053 33201 18117
rect 32985 18031 33201 18053
rect 35758 18127 35923 18147
rect 35758 18068 35784 18127
rect 35896 18068 35923 18127
rect 35758 18043 35923 18068
rect 336 17979 560 18005
rect 441 17675 524 17685
rect 212 17616 301 17621
rect 212 17561 231 17616
rect 284 17561 301 17616
rect 441 17618 451 17675
rect 514 17618 524 17675
rect 441 17608 524 17618
rect 212 17555 301 17561
rect 212 17545 294 17555
rect -1344 17489 294 17545
rect -1344 15921 -1007 17489
rect 2128 17300 2352 17315
rect 2128 17214 2184 17300
rect 2296 17214 2352 17300
rect 2128 17195 2352 17214
rect 6830 17291 7055 17313
rect 6830 17221 6888 17291
rect 7000 17221 7055 17291
rect 6830 17195 7055 17221
rect 11704 17282 11928 17314
rect 11704 17212 11761 17282
rect 11872 17212 11928 17282
rect 11704 17195 11928 17212
rect 16564 17278 16708 17295
rect 16564 17219 16599 17278
rect 16671 17219 16708 17278
rect 16564 17199 16708 17219
rect 21380 17285 21525 17299
rect 21380 17212 21407 17285
rect 21487 17212 21525 17285
rect 21380 17201 21525 17212
rect 26223 17285 26419 17304
rect 26223 17214 26270 17285
rect 26369 17214 26419 17285
rect 26223 17200 26419 17214
rect 31024 17279 31248 17294
rect 31024 17221 31080 17279
rect 31192 17221 31248 17279
rect 31024 17204 31248 17221
rect 37099 17289 37264 17304
rect 37099 17220 37143 17289
rect 37219 17220 37264 17289
rect 37099 17208 37264 17220
rect 2128 16181 2352 16203
rect 2128 16117 2184 16181
rect 2296 16117 2352 16181
rect 2128 16083 2352 16117
rect 6832 16173 7057 16200
rect 6832 16104 6887 16173
rect 7000 16104 7057 16173
rect 6832 16082 7057 16104
rect 11704 16180 11929 16203
rect 11704 16110 11762 16180
rect 11873 16110 11929 16180
rect 11704 16083 11929 16110
rect 16560 16175 16704 16193
rect 16560 16114 16588 16175
rect 16667 16114 16704 16175
rect 16560 16097 16704 16114
rect 21366 16181 21537 16197
rect 21366 16108 21411 16181
rect 21491 16108 21537 16181
rect 21366 16093 21537 16108
rect 26234 16176 26408 16192
rect 26234 16105 26271 16176
rect 26370 16105 26408 16176
rect 26234 16088 26408 16105
rect 31024 16171 31248 16187
rect 31024 16115 31080 16171
rect 31192 16115 31248 16171
rect 31024 16097 31248 16115
rect 37096 16175 37261 16191
rect 37096 16111 37144 16175
rect 37218 16111 37261 16175
rect 37096 16095 37261 16111
rect -1344 15849 512 15921
rect -1344 12051 -1007 15849
rect 440 15793 512 15849
rect 432 15779 519 15793
rect 432 15724 450 15779
rect 505 15724 519 15779
rect 432 15710 519 15724
rect 335 15321 561 15359
rect 335 15254 378 15321
rect 513 15254 561 15321
rect 335 15232 561 15254
rect 3808 15332 4034 15373
rect 3808 15255 3863 15332
rect 3977 15255 4034 15332
rect 3808 15231 4034 15255
rect 8624 15343 8849 15372
rect 8624 15249 8679 15343
rect 8791 15249 8849 15343
rect 8624 15218 8849 15249
rect 13846 15338 14056 15369
rect 13846 15263 13887 15338
rect 14008 15263 14056 15338
rect 13846 15233 14056 15263
rect 18235 15336 18394 15369
rect 18235 15261 18267 15336
rect 18351 15261 18394 15336
rect 18235 15236 18394 15261
rect 23409 15324 23633 15368
rect 23409 15258 23462 15324
rect 23577 15258 23633 15324
rect 23409 15233 23633 15258
rect 27832 15334 28056 15371
rect 27832 15263 27888 15334
rect 28000 15263 28056 15334
rect 27832 15235 28056 15263
rect 32988 15339 33204 15360
rect 32988 15269 33040 15339
rect 33152 15269 33204 15339
rect 32988 15252 33204 15269
rect 35755 15333 35920 15357
rect 35755 15274 35784 15333
rect 35896 15274 35920 15333
rect 35755 15253 35920 15274
rect 210 14821 296 14833
rect 210 14765 224 14821
rect 280 14765 296 14821
rect 210 14750 296 14765
rect 2128 14495 2352 14515
rect 2128 14425 2184 14495
rect 2296 14425 2352 14495
rect 2128 14395 2352 14425
rect 6832 14489 7056 14515
rect 6832 14420 6888 14489
rect 7001 14420 7056 14489
rect 6832 14395 7056 14420
rect 11704 14494 11929 14515
rect 11704 14418 11760 14494
rect 11873 14418 11929 14494
rect 11704 14395 11929 14418
rect 16555 14478 16714 14499
rect 16555 14417 16592 14478
rect 16671 14417 16714 14478
rect 16555 14401 16714 14417
rect 21358 14481 21529 14504
rect 21358 14410 21397 14481
rect 21484 14410 21529 14481
rect 21358 14400 21529 14410
rect 26228 14483 26402 14503
rect 26228 14414 26265 14483
rect 26371 14414 26402 14483
rect 26228 14399 26402 14414
rect 31024 14479 31249 14498
rect 31024 14423 31080 14479
rect 31192 14423 31249 14479
rect 31024 14406 31249 14423
rect 37105 14489 37272 14508
rect 37105 14425 37150 14489
rect 37224 14425 37272 14489
rect 37105 14405 37272 14425
rect 2128 13383 2352 13403
rect 2128 13310 2184 13383
rect 2296 13310 2352 13383
rect 2128 13283 2352 13310
rect 6832 13374 7056 13403
rect 6832 13305 6885 13374
rect 7001 13305 7056 13374
rect 6832 13283 7056 13305
rect 11704 13384 11929 13402
rect 11704 13308 11760 13384
rect 11873 13308 11929 13384
rect 11704 13283 11929 13308
rect 16547 13372 16706 13392
rect 16547 13308 16594 13372
rect 16668 13308 16706 13372
rect 16547 13294 16706 13308
rect 21375 13376 21526 13393
rect 21375 13305 21406 13376
rect 21493 13305 21526 13376
rect 21375 13288 21526 13305
rect 26228 13380 26410 13396
rect 26228 13311 26267 13380
rect 26373 13311 26410 13380
rect 26228 13292 26410 13311
rect 31024 13370 31249 13390
rect 31024 13310 31080 13370
rect 31192 13310 31249 13370
rect 31024 13298 31249 13310
rect 37107 13376 37274 13394
rect 37107 13308 37148 13376
rect 37226 13308 37274 13376
rect 37107 13291 37274 13308
rect 3807 12535 4033 12574
rect 363 12463 532 12498
rect 363 12402 396 12463
rect 501 12402 532 12463
rect 3807 12464 3864 12535
rect 3977 12464 4033 12535
rect 3807 12432 4033 12464
rect 8624 12549 8849 12574
rect 8624 12455 8681 12549
rect 8793 12455 8849 12549
rect 8624 12429 8849 12455
rect 13830 12535 14058 12579
rect 13830 12460 13885 12535
rect 14006 12460 14058 12535
rect 13830 12432 14058 12460
rect 18216 12530 18394 12566
rect 18216 12455 18268 12530
rect 18352 12455 18394 12530
rect 18216 12431 18394 12455
rect 23408 12526 23633 12555
rect 23408 12460 23462 12526
rect 23577 12460 23633 12526
rect 23408 12432 23633 12460
rect 27833 12527 28055 12559
rect 27833 12456 27889 12527
rect 28001 12456 28055 12527
rect 27833 12431 28055 12456
rect 33004 12535 33183 12558
rect 33004 12465 33040 12535
rect 33152 12465 33183 12535
rect 33004 12445 33183 12465
rect 35750 12524 35932 12542
rect 35750 12465 35784 12524
rect 35896 12465 35932 12524
rect 35750 12442 35932 12465
rect 363 12379 532 12402
rect 428 12051 523 12054
rect -1344 12043 523 12051
rect -1344 11987 450 12043
rect 507 11987 523 12043
rect -1344 11983 523 11987
rect -1344 10098 -1007 11983
rect 428 11975 523 11983
rect 2128 11700 2352 11715
rect 2128 11616 2184 11700
rect 2296 11616 2352 11700
rect 2128 11595 2352 11616
rect 6832 11684 7056 11714
rect 6832 11615 6886 11684
rect 7002 11615 7056 11684
rect 6832 11594 7056 11615
rect 11704 11686 11929 11714
rect 11704 11611 11760 11686
rect 11872 11611 11929 11686
rect 11704 11595 11929 11611
rect 16567 11681 16716 11697
rect 16567 11617 16601 11681
rect 16675 11617 16716 11681
rect 16567 11603 16716 11617
rect 21365 11686 21516 11704
rect 21365 11610 21397 11686
rect 21483 11610 21516 11686
rect 21365 11599 21516 11610
rect 26230 11687 26412 11703
rect 26230 11611 26278 11687
rect 26367 11611 26412 11687
rect 26230 11599 26412 11611
rect 31024 11685 31248 11698
rect 31024 11625 31080 11685
rect 31192 11625 31248 11685
rect 31024 11610 31248 11625
rect 37094 11686 37270 11704
rect 37094 11618 37146 11686
rect 37224 11618 37270 11686
rect 37094 11603 37270 11618
rect 31025 10736 31249 10824
rect 2128 10581 2352 10603
rect 2128 10503 2184 10581
rect 2296 10503 2352 10581
rect 2128 10483 2352 10503
rect 6831 10576 7055 10602
rect 6831 10505 6887 10576
rect 7001 10505 7055 10576
rect 6831 10482 7055 10505
rect 11704 10583 11928 10603
rect 11704 10508 11760 10583
rect 11872 10508 11928 10583
rect 11704 10483 11928 10508
rect 16560 10574 16709 10592
rect 16560 10512 16593 10574
rect 16669 10512 16709 10574
rect 16560 10498 16709 10512
rect 21357 10576 21525 10591
rect 21357 10500 21402 10576
rect 21488 10500 21525 10576
rect 21357 10489 21525 10500
rect 26228 10582 26415 10596
rect 26228 10506 26277 10582
rect 26366 10506 26415 10582
rect 26228 10489 26415 10506
rect 31024 10574 31248 10590
rect 31024 10518 31080 10574
rect 31193 10518 31248 10574
rect 31024 10502 31248 10518
rect 37093 10579 37269 10594
rect 37093 10506 37137 10579
rect 37219 10506 37269 10579
rect 37093 10493 37269 10506
rect 447 10178 530 10188
rect 447 10123 461 10178
rect 516 10123 530 10178
rect 447 10115 530 10123
rect 447 10098 524 10115
rect -1344 10026 524 10098
rect -1344 6478 -1007 10026
rect 452 10025 524 10026
rect 336 9719 503 9744
rect 336 9654 368 9719
rect 474 9654 503 9719
rect 336 9632 503 9654
rect 3808 9741 4034 9767
rect 3808 9670 3863 9741
rect 3976 9670 4034 9741
rect 3808 9632 4034 9670
rect 8622 9730 8847 9762
rect 8622 9647 8680 9730
rect 8794 9647 8847 9730
rect 8622 9617 8847 9647
rect 13830 9735 14058 9780
rect 13830 9663 13887 9735
rect 14004 9663 14058 9735
rect 13830 9633 14058 9663
rect 18213 9735 18391 9766
rect 18213 9655 18265 9735
rect 18353 9655 18391 9735
rect 18213 9631 18391 9655
rect 23407 9726 23632 9763
rect 23407 9663 23463 9726
rect 23578 9663 23632 9726
rect 23407 9640 23632 9663
rect 27833 9733 28055 9762
rect 27833 9663 27888 9733
rect 28000 9663 28055 9733
rect 27833 9634 28055 9663
rect 33003 9732 33182 9760
rect 33003 9666 33031 9732
rect 33143 9666 33182 9732
rect 33003 9647 33182 9666
rect 35745 9732 35927 9755
rect 35745 9674 35784 9732
rect 35896 9674 35927 9732
rect 35745 9655 35927 9674
rect 334 9278 419 9288
rect 334 9214 344 9278
rect 408 9214 419 9278
rect 334 9203 419 9214
rect 2128 8893 2352 8915
rect 2128 8813 2184 8893
rect 2296 8813 2352 8893
rect 2128 8795 2352 8813
rect 6833 8885 7057 8913
rect 6833 8814 6886 8885
rect 7000 8814 7057 8885
rect 6833 8795 7057 8814
rect 11704 8889 11928 8914
rect 11704 8811 11760 8889
rect 11872 8811 11928 8889
rect 11704 8794 11928 8811
rect 16551 8878 16727 8900
rect 16551 8816 16598 8878
rect 16674 8816 16727 8878
rect 16551 8802 16727 8816
rect 21357 8885 21525 8904
rect 21357 8811 21397 8885
rect 21484 8811 21525 8885
rect 21357 8802 21525 8811
rect 26223 8886 26410 8907
rect 26223 8811 26265 8886
rect 26364 8811 26410 8886
rect 26223 8800 26410 8811
rect 31033 8882 31231 8900
rect 31033 8826 31079 8882
rect 31192 8826 31231 8882
rect 31033 8807 31231 8826
rect 37092 8885 37270 8901
rect 37092 8812 37142 8885
rect 37224 8812 37270 8885
rect 37092 8802 37270 8812
rect 2128 7784 2352 7803
rect 2128 7714 2184 7784
rect 2296 7714 2352 7784
rect 2128 7683 2352 7714
rect 6832 7773 7056 7802
rect 6832 7708 6888 7773
rect 7000 7708 7056 7773
rect 6832 7684 7056 7708
rect 11704 7781 11928 7802
rect 11704 7703 11760 7781
rect 11872 7703 11928 7781
rect 11704 7683 11928 7703
rect 16540 7772 16716 7791
rect 16540 7706 16589 7772
rect 16670 7706 16716 7772
rect 16540 7693 16716 7706
rect 21363 7779 21532 7793
rect 21363 7705 21404 7779
rect 21491 7705 21532 7779
rect 21363 7689 21532 7705
rect 26231 7783 26414 7796
rect 26231 7708 26273 7783
rect 26372 7708 26414 7783
rect 26231 7693 26414 7708
rect 31031 7772 31229 7790
rect 31031 7716 31079 7772
rect 31192 7716 31229 7772
rect 31031 7697 31229 7716
rect 37097 7779 37275 7794
rect 37097 7711 37144 7779
rect 37228 7711 37275 7779
rect 37097 7695 37275 7711
rect 3807 6935 4033 6967
rect 337 6874 561 6900
rect 337 6805 390 6874
rect 505 6805 561 6874
rect 3807 6854 3863 6935
rect 3977 6854 4033 6935
rect 3807 6832 4033 6854
rect 8623 6928 8848 6965
rect 8623 6849 8679 6928
rect 8791 6849 8848 6928
rect 8623 6824 8848 6849
rect 13832 6938 14058 6973
rect 13832 6866 13886 6938
rect 14003 6866 14058 6938
rect 13832 6838 14058 6866
rect 18225 6956 18392 6977
rect 18225 6876 18263 6956
rect 18351 6876 18392 6956
rect 18225 6855 18392 6876
rect 23406 6928 23634 6962
rect 23406 6865 23462 6928
rect 23577 6865 23634 6928
rect 23406 6834 23634 6865
rect 27831 6939 28053 6967
rect 27831 6869 27887 6939
rect 27999 6869 28053 6939
rect 27831 6832 28053 6869
rect 33009 6930 33190 6951
rect 33009 6864 33041 6930
rect 33153 6864 33190 6930
rect 33009 6842 33190 6864
rect 35737 6921 35937 6945
rect 35737 6863 35784 6921
rect 35896 6863 35937 6921
rect 35737 6839 35937 6863
rect 337 6779 561 6805
rect 320 6478 406 6482
rect -1344 6473 406 6478
rect -1344 6421 334 6473
rect 389 6421 406 6473
rect -1344 6415 406 6421
rect -1344 4735 -1007 6415
rect 320 6408 406 6415
rect 544 6479 628 6489
rect 544 6416 554 6479
rect 618 6416 628 6479
rect 544 6406 628 6416
rect 2128 6088 2352 6115
rect 2128 6012 2184 6088
rect 2296 6012 2352 6088
rect 2128 5995 2352 6012
rect 6832 6081 7056 6115
rect 6832 6016 6888 6081
rect 7000 6016 7056 6081
rect 6832 5995 7056 6016
rect 11703 6089 11927 6114
rect 11703 6016 11761 6089
rect 11874 6016 11927 6089
rect 11703 5995 11927 6016
rect 16558 6082 16730 6104
rect 16558 6016 16593 6082
rect 16674 6016 16730 6082
rect 16558 5998 16730 6016
rect 21359 6083 21528 6105
rect 21359 6011 21400 6083
rect 21485 6011 21528 6083
rect 21359 6001 21528 6011
rect 26232 6090 26415 6102
rect 26232 6010 26275 6090
rect 26367 6010 26415 6090
rect 26232 5999 26415 6010
rect 31049 6082 31220 6098
rect 31049 6026 31080 6082
rect 31193 6026 31220 6082
rect 31049 6009 31220 6026
rect 37090 6083 37270 6101
rect 37090 6015 37140 6083
rect 37224 6015 37270 6083
rect 37090 6002 37270 6015
rect 2128 4984 2353 5003
rect 2128 4910 2184 4984
rect 2296 4910 2353 4984
rect 2128 4883 2353 4910
rect 6832 4974 7056 5003
rect 6832 4903 6888 4974
rect 7001 4903 7056 4974
rect 6832 4883 7056 4903
rect 11704 4980 11929 5002
rect 11704 4907 11759 4980
rect 11872 4907 11929 4980
rect 11704 4883 11929 4907
rect 16545 4976 16717 4993
rect 16545 4906 16589 4976
rect 16672 4906 16717 4976
rect 16545 4887 16717 4906
rect 21375 4974 21532 4993
rect 21375 4902 21408 4974
rect 21493 4902 21532 4974
rect 21375 4887 21532 4902
rect 26242 4980 26415 4996
rect 26242 4900 26281 4980
rect 26373 4900 26415 4980
rect 31050 4977 31221 4990
rect 31050 4921 31080 4977
rect 31192 4921 31221 4977
rect 31050 4901 31221 4921
rect 37100 4976 37280 4992
rect 37100 4910 37140 4976
rect 37228 4910 37280 4976
rect 26242 4886 26415 4900
rect 37100 4893 37280 4910
rect -1344 4663 618 4735
rect -1344 2800 -1007 4663
rect 546 4590 618 4663
rect 536 4577 626 4590
rect 536 4523 557 4577
rect 611 4523 626 4577
rect 536 4506 626 4523
rect 336 4141 561 4200
rect 336 4062 390 4141
rect 507 4062 561 4141
rect 336 4028 561 4062
rect 3808 4139 4032 4172
rect 3808 4058 3863 4139
rect 3977 4058 4032 4139
rect 3808 4031 4032 4058
rect 8624 4129 8849 4164
rect 8624 4052 8680 4129
rect 8793 4052 8849 4129
rect 8624 4025 8849 4052
rect 13831 4135 14057 4166
rect 13831 4060 13887 4135
rect 14000 4060 14057 4135
rect 13831 4033 14057 4060
rect 18222 4141 18389 4170
rect 18222 4066 18267 4141
rect 18360 4066 18389 4141
rect 18222 4048 18389 4066
rect 23407 4127 23635 4161
rect 23407 4056 23460 4127
rect 23576 4056 23635 4127
rect 23407 4033 23635 4056
rect 27834 4123 28056 4160
rect 27834 4050 27887 4123
rect 28001 4050 28056 4123
rect 27834 4025 28056 4050
rect 32997 4136 33178 4158
rect 32997 4072 33030 4136
rect 33139 4072 33178 4136
rect 32997 4049 33178 4072
rect 35742 4130 35942 4159
rect 35742 4074 35783 4130
rect 35896 4074 35942 4130
rect 35742 4053 35942 4074
rect 318 3677 401 3687
rect 318 3617 328 3677
rect 391 3617 401 3677
rect 318 3607 401 3617
rect 2128 3293 2352 3315
rect 2128 3214 2184 3293
rect 2296 3214 2352 3293
rect 2128 3195 2352 3214
rect 6832 3288 7056 3314
rect 6832 3217 6888 3288
rect 7001 3217 7056 3288
rect 6832 3194 7056 3217
rect 11701 3284 11926 3314
rect 11701 3209 11757 3284
rect 11875 3209 11926 3284
rect 11701 3195 11926 3209
rect 16560 3288 16719 3302
rect 16560 3218 16594 3288
rect 16677 3218 16719 3288
rect 16560 3202 16719 3218
rect 21371 3283 21528 3303
rect 21371 3212 21401 3283
rect 21486 3212 21528 3283
rect 21371 3197 21528 3212
rect 26229 3290 26402 3309
rect 26229 3210 26264 3290
rect 26360 3210 26402 3290
rect 26229 3199 26402 3210
rect 31051 3278 31233 3299
rect 31051 3222 31080 3278
rect 31192 3222 31233 3278
rect 31051 3204 31233 3222
rect 37093 3285 37278 3305
rect 37093 3219 37137 3285
rect 37225 3219 37278 3285
rect 37093 3206 37278 3219
rect 2128 2172 2352 2203
rect 2128 2104 2184 2172
rect 2296 2104 2352 2172
rect 2128 2083 2352 2104
rect 6832 2173 7056 2204
rect 6832 2104 6887 2173
rect 7001 2104 7056 2173
rect 6832 2084 7056 2104
rect 11702 2181 11929 2200
rect 11702 2106 11758 2181
rect 11876 2106 11929 2181
rect 11702 2085 11929 2106
rect 16553 2177 16712 2194
rect 16553 2104 16595 2177
rect 16675 2104 16712 2177
rect 16553 2094 16712 2104
rect 21376 2174 21524 2196
rect 21376 2103 21403 2174
rect 21488 2103 21524 2174
rect 21376 2084 21524 2103
rect 26227 2179 26412 2195
rect 26227 2099 26276 2179
rect 26372 2099 26412 2179
rect 31046 2178 31228 2194
rect 31046 2117 31079 2178
rect 31193 2117 31228 2178
rect 31046 2099 31228 2117
rect 26227 2088 26412 2099
rect 3808 1332 4032 1378
rect 3808 1265 3864 1332
rect 3976 1265 4032 1332
rect 3808 1232 4032 1265
rect 8625 1334 8849 1364
rect 8625 1257 8679 1334
rect 8792 1257 8849 1334
rect 8625 1231 8849 1257
rect 13834 1328 14055 1363
rect 13834 1255 13872 1328
rect 14002 1255 14055 1328
rect 13834 1219 14055 1255
rect 18198 1335 18424 1361
rect 18198 1260 18262 1335
rect 18355 1260 18424 1335
rect 18198 1233 18424 1260
rect 23409 1342 23632 1368
rect 23409 1271 23462 1342
rect 23578 1271 23632 1342
rect 23409 1233 23632 1271
rect 27832 1330 28059 1357
rect 27832 1257 27887 1330
rect 28001 1257 28059 1330
rect 27832 1233 28059 1257
rect 33008 1329 33186 1356
rect 33008 1265 33043 1329
rect 33152 1265 33186 1329
rect 33008 1241 33186 1265
rect 2128 489 2352 515
rect 2128 416 2184 489
rect 2296 416 2352 489
rect 2128 395 2352 416
rect 6831 487 7057 515
rect 6831 418 6887 487
rect 7001 418 7057 487
rect 6831 395 7057 418
rect 11704 487 11931 511
rect 11704 410 11760 487
rect 11872 410 11931 487
rect 11704 396 11931 410
rect 16529 485 16723 502
rect 16529 412 16588 485
rect 16668 412 16723 485
rect 16529 401 16723 412
rect 21369 480 21517 507
rect 21369 408 21402 480
rect 21481 408 21517 480
rect 21369 395 21517 408
rect 26229 483 26414 505
rect 26229 406 26275 483
rect 26363 406 26414 483
rect 26229 398 26414 406
rect 31041 482 31228 504
rect 31041 421 31079 482
rect 31193 421 31228 482
rect 31041 402 31228 421
<< via2 >>
rect 3528 26656 3640 26767
rect 17300 26600 17418 26707
rect 35784 27796 35874 27869
rect 35801 26846 35890 26918
rect 35794 25881 35883 25953
rect 35800 24915 35893 24993
rect 40384 29049 40502 29131
rect 37124 27023 37213 27079
rect 37123 26063 37244 26128
rect 37126 25104 37244 25163
rect 472 24324 530 24380
rect 391 22657 504 22733
rect 3881 22614 3971 22672
rect 8680 23169 8793 23243
rect 13888 23184 13944 23240
rect 10358 22848 10418 22850
rect 10358 22794 10361 22848
rect 10361 22794 10415 22848
rect 10415 22794 10418 22848
rect 10358 22792 10418 22794
rect 18283 23184 18339 23240
rect 20104 24360 20160 24416
rect 23493 23184 23549 23240
rect 25144 24360 25200 24416
rect 27862 23179 28000 23251
rect 37119 24130 37237 24189
rect 29788 22792 29852 22852
rect 11761 22389 11874 22465
rect 16605 22400 16661 22456
rect 21421 22400 21477 22456
rect 26292 22400 26348 22456
rect 31111 22400 31167 22456
rect 3862 22224 3923 22226
rect 3862 22172 3865 22224
rect 3865 22172 3920 22224
rect 3920 22172 3923 22224
rect 3862 22170 3923 22172
rect 2184 21703 2296 21777
rect 6887 21698 7001 21776
rect 11760 21700 11873 21782
rect 16593 21710 16683 21769
rect 21412 21709 21490 21773
rect 26264 21706 26375 21776
rect 31080 21714 31193 21771
rect 37146 21707 37224 21773
rect 467 21377 528 21380
rect 467 21325 470 21377
rect 470 21325 525 21377
rect 525 21325 528 21377
rect 467 21323 528 21325
rect 392 20849 505 20925
rect 3864 20871 3976 20940
rect 8678 20855 8793 20940
rect 13889 20866 14003 20934
rect 18268 20864 18348 20943
rect 23462 20862 23576 20944
rect 27887 20864 28000 20937
rect 33039 20874 33155 20938
rect 35784 20869 35896 20928
rect 2184 20019 2296 20085
rect 6888 20014 7000 20091
rect 11760 20016 11872 20098
rect 16583 20022 16673 20081
rect 21409 20021 21486 20085
rect 26277 20017 26366 20089
rect 31079 20020 31192 20077
rect 37145 20023 37223 20089
rect 2184 18907 2296 18973
rect 6888 18901 7000 18976
rect 11760 18904 11872 18986
rect 16593 18910 16665 18969
rect 21404 18914 21481 18978
rect 26281 18903 26370 18975
rect 31080 18911 31192 18969
rect 37151 18909 37227 18978
rect 392 18005 505 18072
rect 3863 18059 3977 18136
rect 8680 18055 8792 18139
rect 13888 18070 14002 18138
rect 18269 18065 18349 18144
rect 23464 18068 23575 18143
rect 27889 18066 28002 18139
rect 33038 18053 33154 18117
rect 35784 18068 35896 18127
rect 451 17673 514 17675
rect 451 17621 454 17673
rect 454 17621 510 17673
rect 510 17621 514 17673
rect 451 17618 514 17621
rect 2184 17214 2296 17300
rect 6888 17221 7000 17291
rect 11761 17212 11872 17282
rect 16599 17219 16671 17278
rect 21407 17212 21487 17285
rect 26270 17214 26369 17285
rect 31080 17221 31192 17279
rect 37143 17220 37219 17289
rect 2184 16117 2296 16181
rect 6887 16104 7000 16173
rect 11762 16110 11873 16180
rect 16588 16114 16667 16175
rect 21411 16108 21491 16181
rect 26271 16105 26370 16176
rect 31080 16115 31192 16171
rect 37144 16111 37218 16175
rect 378 15254 513 15321
rect 3863 15255 3977 15332
rect 8679 15249 8791 15343
rect 13887 15263 14008 15338
rect 18267 15261 18351 15336
rect 23462 15258 23577 15324
rect 27888 15263 28000 15334
rect 33040 15269 33152 15339
rect 35784 15274 35896 15333
rect 224 14819 280 14821
rect 224 14765 280 14819
rect 2184 14425 2296 14495
rect 6888 14420 7001 14489
rect 11760 14418 11873 14494
rect 16592 14417 16671 14478
rect 21397 14410 21484 14481
rect 26265 14414 26371 14483
rect 31080 14423 31192 14479
rect 37150 14425 37224 14489
rect 2184 13310 2296 13383
rect 6885 13305 7001 13374
rect 11760 13308 11873 13384
rect 16594 13308 16668 13372
rect 21406 13305 21493 13376
rect 26267 13311 26373 13380
rect 31080 13310 31192 13370
rect 37148 13308 37226 13376
rect 396 12402 501 12463
rect 3864 12464 3977 12535
rect 8681 12455 8793 12549
rect 13885 12460 14006 12535
rect 18268 12455 18352 12530
rect 23462 12460 23577 12526
rect 27889 12456 28001 12527
rect 33040 12465 33152 12535
rect 35784 12465 35896 12524
rect 2184 11616 2296 11700
rect 6886 11615 7002 11684
rect 11760 11611 11872 11686
rect 16601 11617 16675 11681
rect 21397 11610 21483 11686
rect 26278 11611 26367 11687
rect 31080 11625 31192 11685
rect 37146 11618 37224 11686
rect 2184 10503 2296 10581
rect 6887 10505 7001 10576
rect 11760 10508 11872 10583
rect 16593 10512 16669 10574
rect 21402 10500 21488 10576
rect 26277 10506 26366 10582
rect 31080 10573 31193 10574
rect 31080 10518 31193 10573
rect 37137 10506 37219 10579
rect 368 9654 474 9719
rect 3863 9670 3976 9741
rect 8680 9647 8794 9730
rect 13887 9663 14004 9735
rect 18265 9655 18353 9735
rect 23463 9663 23578 9726
rect 27888 9663 28000 9733
rect 33031 9666 33143 9732
rect 35784 9674 35896 9732
rect 344 9274 408 9278
rect 344 9217 347 9274
rect 347 9217 404 9274
rect 404 9217 408 9274
rect 344 9214 408 9217
rect 2184 8813 2296 8893
rect 6886 8814 7000 8885
rect 11760 8811 11872 8889
rect 16598 8816 16674 8878
rect 21397 8811 21484 8885
rect 26265 8811 26364 8886
rect 31079 8826 31192 8882
rect 37142 8812 37224 8885
rect 2184 7714 2296 7784
rect 6888 7708 7000 7773
rect 11760 7703 11872 7781
rect 16589 7706 16670 7772
rect 21404 7705 21491 7779
rect 26273 7708 26372 7783
rect 31079 7716 31192 7772
rect 37144 7711 37228 7779
rect 390 6805 505 6874
rect 3863 6854 3977 6935
rect 8679 6849 8791 6928
rect 13886 6866 14003 6938
rect 18263 6876 18351 6956
rect 23462 6865 23577 6928
rect 27887 6869 27999 6939
rect 33041 6864 33153 6930
rect 35784 6863 35896 6921
rect 554 6416 618 6479
rect 2184 6012 2296 6088
rect 6888 6016 7000 6081
rect 11761 6016 11874 6089
rect 16593 6016 16674 6082
rect 21400 6011 21485 6083
rect 26275 6010 26367 6090
rect 31080 6026 31193 6082
rect 37140 6015 37224 6083
rect 2184 4910 2296 4984
rect 6888 4903 7001 4974
rect 11759 4907 11872 4980
rect 16589 4906 16672 4976
rect 21408 4902 21493 4974
rect 26281 4900 26373 4980
rect 31080 4921 31192 4977
rect 37140 4910 37228 4976
rect 390 4062 507 4141
rect 3863 4058 3977 4139
rect 8680 4052 8793 4129
rect 13887 4060 14000 4135
rect 18267 4066 18360 4141
rect 23460 4056 23576 4127
rect 27887 4050 28001 4123
rect 33030 4072 33139 4136
rect 35783 4074 35896 4130
rect 328 3674 391 3677
rect 328 3620 333 3674
rect 333 3620 388 3674
rect 388 3620 391 3674
rect 328 3617 391 3620
rect 2184 3214 2296 3293
rect 6888 3217 7001 3288
rect 11757 3209 11875 3284
rect 16594 3218 16677 3288
rect 21401 3212 21486 3283
rect 26264 3210 26360 3290
rect 31080 3222 31192 3278
rect 37137 3219 37225 3285
rect 2184 2104 2296 2172
rect 6887 2104 7001 2173
rect 11758 2106 11876 2181
rect 16595 2104 16675 2177
rect 21403 2103 21488 2174
rect 26276 2099 26372 2179
rect 31079 2117 31193 2178
rect 3864 1265 3976 1332
rect 8679 1257 8792 1334
rect 13872 1255 14002 1328
rect 18262 1260 18355 1335
rect 23462 1271 23578 1342
rect 27887 1257 28001 1330
rect 33043 1265 33152 1329
rect 2184 416 2296 489
rect 6887 418 7001 487
rect 11760 410 11872 487
rect 16588 412 16668 485
rect 21402 408 21481 480
rect 26275 406 26363 483
rect 31079 421 31193 482
<< metal3 >>
rect -10148 36995 -7674 37008
rect 48434 36995 50908 37079
rect -10148 34395 50919 36995
rect -10148 18432 -7674 34395
rect 2071 28125 2408 34395
rect 2071 27854 2120 28125
rect 2373 27854 2408 28125
rect 2071 27782 2408 27854
rect 6805 27952 7142 34395
rect 6805 27707 6889 27952
rect 7064 27707 7142 27952
rect 11652 28436 11989 34395
rect 11652 28067 11691 28436
rect 11959 28067 11989 28436
rect 11652 27734 11989 28067
rect 16465 28508 16802 34395
rect 16465 28225 16525 28508
rect 16765 28225 16802 28508
rect 16465 28021 16802 28225
rect 21284 28583 21621 34395
rect 21284 28222 21331 28583
rect 21592 28222 21621 28583
rect 21284 28111 21621 28222
rect 26158 28269 26495 34395
rect 26158 27940 26205 28269
rect 26457 27940 26495 28269
rect 6805 27579 7142 27707
rect 26158 27671 26495 27940
rect 30980 28484 31317 34395
rect 30980 28204 31016 28484
rect 31278 28204 31317 28484
rect 30980 27930 31317 28204
rect 35755 27869 35905 27885
rect 35755 27796 35784 27869
rect 35874 27796 35905 27869
rect 35755 27786 35905 27796
rect 37007 27079 37344 34395
rect 40321 29131 40543 29198
rect 40321 29049 40384 29131
rect 40502 29049 40543 29131
rect 40321 28997 40543 29049
rect 37007 27023 37124 27079
rect 37213 27023 37344 27079
rect 35768 26918 35918 26931
rect 35768 26846 35801 26918
rect 35890 26846 35918 26918
rect 35768 26832 35918 26846
rect 3414 26824 3761 26825
rect -1736 26767 3761 26824
rect -1736 26656 3528 26767
rect 3640 26656 3761 26767
rect -1736 26600 3761 26656
rect 17191 26707 17530 26769
rect 17191 26600 17300 26707
rect 17418 26600 17530 26707
rect 37007 26694 37344 27023
rect -1736 25396 -1400 26600
rect 17191 26487 17530 26600
rect -1736 21384 -1399 25396
rect 6473 24585 7469 24588
rect 17248 24585 17472 26487
rect 37106 26128 37262 26143
rect 37106 26063 37123 26128
rect 37244 26063 37262 26128
rect 37106 26050 37262 26063
rect 35772 25953 35906 25968
rect 35772 25881 35794 25953
rect 35883 25881 35906 25953
rect 35772 25873 35906 25881
rect 37106 25163 37262 25179
rect 37106 25104 37126 25163
rect 37244 25104 37262 25163
rect 37106 25086 37262 25104
rect 35790 24993 35903 25003
rect 35790 24915 35800 24993
rect 35893 24915 35903 24993
rect 35790 24905 35903 24915
rect 224 24416 30070 24585
rect 224 24380 20104 24416
rect 224 24324 472 24380
rect 530 24360 20104 24380
rect 20160 24360 25144 24416
rect 25200 24360 30070 24416
rect 530 24324 30070 24360
rect 224 24248 30070 24324
rect 2022 24247 2541 24248
rect 336 22733 562 22762
rect 336 22657 391 22733
rect 504 22657 562 22733
rect 336 22628 562 22657
rect 3633 22237 3710 24248
rect 8624 23243 8847 23275
rect 8624 23169 8680 23243
rect 8793 23169 8847 23243
rect 8624 23154 8847 23169
rect 10352 22860 10424 24248
rect 11310 24247 12106 24248
rect 16409 24247 16979 24248
rect 27843 23251 28014 23274
rect 13878 23240 13954 23250
rect 13878 23184 13888 23240
rect 13944 23184 13954 23240
rect 13878 23174 13954 23184
rect 18273 23240 18349 23250
rect 18273 23184 18283 23240
rect 18339 23184 18349 23240
rect 18273 23174 18349 23184
rect 23483 23240 23559 23250
rect 23483 23184 23493 23240
rect 23549 23184 23559 23240
rect 23483 23174 23559 23184
rect 27843 23179 27862 23251
rect 28000 23179 28014 23251
rect 27843 23158 28014 23179
rect 29782 22862 29854 24248
rect 37086 24189 37271 24207
rect 37086 24130 37119 24189
rect 37237 24130 37271 24189
rect 37086 24118 37271 24130
rect 10348 22850 10428 22860
rect 10348 22792 10358 22850
rect 10418 22792 10428 22850
rect 10348 22782 10428 22792
rect 29778 22852 29862 22862
rect 29778 22792 29788 22852
rect 29852 22792 29862 22852
rect 29778 22782 29862 22792
rect 3836 22672 4021 22707
rect 3836 22614 3881 22672
rect 3971 22614 4021 22672
rect 3836 22586 4021 22614
rect 11727 22465 11904 22491
rect 11727 22389 11761 22465
rect 11874 22389 11904 22465
rect 16595 22456 16671 22466
rect 16595 22400 16605 22456
rect 16661 22400 16671 22456
rect 16595 22390 16671 22400
rect 21411 22456 21487 22466
rect 21411 22400 21421 22456
rect 21477 22400 21487 22456
rect 21411 22390 21487 22400
rect 26282 22456 26358 22466
rect 26282 22400 26292 22456
rect 26348 22400 26358 22456
rect 26282 22390 26358 22400
rect 31101 22456 31177 22466
rect 31101 22400 31111 22456
rect 31167 22400 31177 22456
rect 31101 22390 31177 22400
rect 11727 22369 11904 22389
rect 3633 22226 3934 22237
rect 3633 22170 3862 22226
rect 3923 22170 3934 22226
rect 3633 22160 3934 22170
rect 3851 22159 3934 22160
rect 2128 21777 2352 21803
rect 2128 21703 2184 21777
rect 2296 21703 2352 21777
rect 2128 21683 2352 21703
rect 6832 21776 7056 21803
rect 6832 21698 6887 21776
rect 7001 21698 7056 21776
rect 6832 21683 7056 21698
rect 11704 21782 11928 21803
rect 11704 21700 11760 21782
rect 11873 21700 11928 21782
rect 11704 21683 11928 21700
rect 16520 21769 16744 21803
rect 16520 21710 16593 21769
rect 16683 21710 16744 21769
rect 16520 21683 16744 21710
rect 21358 21773 21543 21792
rect 21358 21709 21412 21773
rect 21490 21709 21543 21773
rect 21358 21696 21543 21709
rect 26222 21776 26412 21792
rect 26222 21706 26264 21776
rect 26375 21706 26412 21776
rect 26222 21687 26412 21706
rect 31024 21771 31248 21792
rect 31024 21714 31080 21771
rect 31193 21714 31248 21771
rect 31024 21691 31248 21714
rect 37107 21773 37270 21793
rect 37107 21707 37146 21773
rect 37224 21707 37270 21773
rect 37107 21692 37270 21707
rect 457 21384 538 21390
rect -1736 21380 538 21384
rect -1736 21323 467 21380
rect 528 21323 538 21380
rect -1736 21317 538 21323
rect -10148 18392 -2944 18432
rect -10148 18260 -3218 18392
rect -3023 18260 -2944 18392
rect -10148 18234 -2944 18260
rect -10148 12867 -7674 18234
rect -1736 17684 -1399 21317
rect 457 21313 538 21317
rect 45018 21224 46209 21546
rect -504 21185 46209 21224
rect -504 21181 27903 21185
rect -504 21105 402 21181
rect 487 21179 27903 21181
rect 487 21105 3887 21179
rect -504 21103 3887 21105
rect 3972 21103 8706 21179
rect 8791 21173 18269 21179
rect 8791 21103 13893 21173
rect -504 21097 13893 21103
rect 13978 21103 18269 21173
rect 18354 21173 27903 21179
rect 18354 21103 23473 21173
rect 13978 21097 23473 21103
rect 23558 21109 27903 21173
rect 27988 21175 46209 21185
rect 27988 21173 35797 21175
rect 27988 21109 33024 21173
rect 23558 21097 33024 21109
rect 33109 21099 35797 21173
rect 35882 21099 46209 21175
rect 33109 21097 46209 21099
rect -504 21056 46209 21097
rect 335 20925 559 20947
rect 335 20849 392 20925
rect 505 20849 559 20925
rect 335 20829 559 20849
rect 3808 20940 4034 20970
rect 3808 20871 3864 20940
rect 3976 20871 4034 20940
rect 3808 20844 4034 20871
rect 8623 20940 8848 20987
rect 8623 20855 8678 20940
rect 8793 20855 8848 20940
rect 8623 20822 8848 20855
rect 13856 20934 14035 20958
rect 13856 20866 13889 20934
rect 14003 20866 14035 20934
rect 13856 20835 14035 20866
rect 18231 20943 18383 20974
rect 18231 20864 18268 20943
rect 18348 20864 18383 20943
rect 18231 20834 18383 20864
rect 23408 20944 23632 20973
rect 23408 20862 23462 20944
rect 23576 20862 23632 20944
rect 23408 20832 23632 20862
rect 27831 20937 28057 20949
rect 27831 20864 27887 20937
rect 28000 20864 28057 20937
rect 27831 20833 28057 20864
rect 32984 20938 33208 20974
rect 32984 20874 33039 20938
rect 33155 20874 33208 20938
rect 32984 20848 33208 20874
rect 35736 20928 35937 20948
rect 35736 20869 35784 20928
rect 35896 20869 35937 20928
rect 35736 20845 35937 20869
rect 45018 20796 46209 21056
rect 2128 20085 2352 20115
rect 2128 20019 2184 20085
rect 2296 20019 2352 20085
rect 2128 19995 2352 20019
rect 6832 20091 7057 20115
rect 6832 20014 6888 20091
rect 7000 20014 7057 20091
rect 6832 19995 7057 20014
rect 11704 20098 11928 20115
rect 11704 20016 11760 20098
rect 11872 20016 11928 20098
rect 11704 19995 11928 20016
rect 16540 20081 16720 20096
rect 16540 20022 16583 20081
rect 16673 20022 16720 20081
rect 16540 20004 16720 20022
rect 21355 20085 21540 20098
rect 21355 20021 21409 20085
rect 21486 20021 21540 20085
rect 21355 20006 21540 20021
rect 26228 20089 26418 20104
rect 26228 20017 26277 20089
rect 26366 20017 26418 20089
rect 26228 19999 26418 20017
rect 31023 20077 31248 20097
rect 31023 20020 31079 20077
rect 31192 20020 31248 20077
rect 31023 20003 31248 20020
rect 37092 20089 37277 20108
rect 37092 20023 37145 20089
rect 37223 20023 37277 20089
rect 37092 20006 37277 20023
rect 2128 18973 2352 19003
rect 2128 18907 2184 18973
rect 2296 18907 2352 18973
rect 2128 18883 2352 18907
rect 6832 18976 7056 19002
rect 6832 18901 6888 18976
rect 7000 18901 7056 18976
rect 6832 18883 7056 18901
rect 11704 18986 11928 19002
rect 11704 18904 11760 18986
rect 11872 18904 11928 18986
rect 11704 18883 11928 18904
rect 16540 18969 16720 18988
rect 16540 18910 16593 18969
rect 16665 18910 16720 18969
rect 16540 18896 16720 18910
rect 21371 18978 21516 18995
rect 21371 18914 21404 18978
rect 21481 18914 21516 18978
rect 21371 18897 21516 18914
rect 26221 18975 26417 18991
rect 26221 18903 26281 18975
rect 26370 18903 26417 18975
rect 26221 18887 26417 18903
rect 31024 18969 31249 18988
rect 31024 18911 31080 18969
rect 31192 18911 31249 18969
rect 31024 18894 31249 18911
rect 37099 18978 37284 18996
rect 37099 18909 37151 18978
rect 37227 18909 37284 18978
rect 37099 18894 37284 18909
rect 48434 18405 50908 34395
rect 45275 18401 50908 18405
rect -322 18382 50908 18401
rect -322 18380 21374 18382
rect -322 18374 11718 18380
rect -322 18368 6871 18374
rect -322 18265 -217 18368
rect -32 18265 2155 18368
rect -322 18258 2155 18265
rect 2326 18264 6871 18368
rect 7042 18270 11718 18374
rect 11889 18368 21374 18380
rect 11889 18270 16548 18368
rect 7042 18264 16548 18270
rect 2326 18258 16548 18264
rect 16719 18262 21374 18368
rect 21545 18378 50908 18382
rect 21545 18374 31048 18378
rect 21545 18262 26231 18374
rect 16719 18258 26231 18262
rect -322 18254 26231 18258
rect 26402 18258 31048 18374
rect 31219 18374 50908 18378
rect 31219 18258 37093 18374
rect 26402 18254 37093 18258
rect 37264 18254 50908 18374
rect -322 18233 50908 18254
rect 3807 18136 4033 18157
rect 336 18072 560 18097
rect 336 18005 392 18072
rect 505 18005 560 18072
rect 3807 18059 3863 18136
rect 3977 18059 4033 18136
rect 3807 18031 4033 18059
rect 8625 18139 8848 18176
rect 8625 18055 8680 18139
rect 8792 18055 8848 18139
rect 8625 18028 8848 18055
rect 13840 18138 14050 18175
rect 13840 18070 13888 18138
rect 14002 18070 14050 18138
rect 13840 18039 14050 18070
rect 18228 18144 18387 18174
rect 18228 18065 18269 18144
rect 18349 18065 18387 18144
rect 18228 18041 18387 18065
rect 23408 18143 23632 18167
rect 23408 18068 23464 18143
rect 23575 18068 23632 18143
rect 23408 18032 23632 18068
rect 27833 18139 28057 18167
rect 27833 18066 27889 18139
rect 28002 18066 28057 18139
rect 27833 18031 28057 18066
rect 32985 18117 33201 18139
rect 32985 18053 33038 18117
rect 33154 18053 33201 18117
rect 32985 18031 33201 18053
rect 35758 18127 35923 18147
rect 35758 18068 35784 18127
rect 35896 18068 35923 18127
rect 35758 18043 35923 18068
rect 336 17979 560 18005
rect 441 17684 524 17685
rect -1736 17675 524 17684
rect -1736 17618 451 17675
rect 514 17618 524 17675
rect -1736 17616 524 17618
rect -1736 14825 -1399 17616
rect 441 17608 524 17616
rect 2128 17300 2352 17315
rect 2128 17214 2184 17300
rect 2296 17214 2352 17300
rect 2128 17195 2352 17214
rect 6830 17291 7055 17313
rect 6830 17221 6888 17291
rect 7000 17221 7055 17291
rect 6830 17195 7055 17221
rect 11704 17282 11928 17314
rect 11704 17212 11761 17282
rect 11872 17212 11928 17282
rect 11704 17195 11928 17212
rect 16564 17278 16708 17295
rect 16564 17219 16599 17278
rect 16671 17219 16708 17278
rect 16564 17199 16708 17219
rect 21380 17285 21525 17299
rect 21380 17212 21407 17285
rect 21487 17212 21525 17285
rect 21380 17201 21525 17212
rect 26223 17285 26419 17304
rect 26223 17214 26270 17285
rect 26369 17214 26419 17285
rect 26223 17200 26419 17214
rect 31024 17279 31248 17294
rect 31024 17221 31080 17279
rect 31192 17221 31248 17279
rect 31024 17204 31248 17221
rect 37099 17289 37264 17304
rect 37099 17220 37143 17289
rect 37219 17220 37264 17289
rect 37099 17208 37264 17220
rect 2128 16181 2352 16203
rect 2128 16117 2184 16181
rect 2296 16117 2352 16181
rect 2128 16083 2352 16117
rect 6832 16173 7057 16200
rect 6832 16104 6887 16173
rect 7000 16104 7057 16173
rect 6832 16082 7057 16104
rect 11704 16180 11929 16203
rect 11704 16110 11762 16180
rect 11873 16110 11929 16180
rect 11704 16083 11929 16110
rect 16560 16175 16704 16193
rect 16560 16114 16588 16175
rect 16667 16114 16704 16175
rect 16560 16097 16704 16114
rect 21366 16181 21537 16197
rect 21366 16108 21411 16181
rect 21491 16108 21537 16181
rect 21366 16093 21537 16108
rect 26234 16176 26408 16192
rect 26234 16105 26271 16176
rect 26370 16105 26408 16176
rect 26234 16088 26408 16105
rect 31024 16171 31248 16187
rect 31024 16115 31080 16171
rect 31192 16115 31248 16171
rect 31024 16097 31248 16115
rect 37096 16175 37261 16191
rect 37096 16111 37144 16175
rect 37218 16111 37261 16175
rect 37096 16095 37261 16111
rect 45014 15653 46079 15924
rect -390 15608 46079 15653
rect -390 15605 35802 15608
rect -390 15603 33057 15605
rect -390 15539 439 15603
rect 503 15600 33057 15603
rect 503 15598 27903 15600
rect 503 15593 18260 15598
rect 503 15539 3877 15593
rect -390 15529 3877 15539
rect 3941 15529 8694 15593
rect 8758 15529 13902 15593
rect 13966 15534 18260 15593
rect 18324 15534 23473 15598
rect 23537 15536 27903 15598
rect 27967 15541 33057 15600
rect 33121 15544 35802 15605
rect 35866 15544 46079 15608
rect 33121 15541 46079 15544
rect 27967 15536 46079 15541
rect 23537 15534 46079 15536
rect 13966 15529 46079 15534
rect -390 15485 46079 15529
rect 335 15321 561 15359
rect 335 15254 378 15321
rect 513 15254 561 15321
rect 335 15232 561 15254
rect 3808 15332 4034 15373
rect 3808 15255 3863 15332
rect 3977 15255 4034 15332
rect 3808 15231 4034 15255
rect 8624 15343 8849 15372
rect 8624 15249 8679 15343
rect 8791 15249 8849 15343
rect 8624 15218 8849 15249
rect 13846 15338 14056 15369
rect 13846 15263 13887 15338
rect 14008 15263 14056 15338
rect 13846 15233 14056 15263
rect 18235 15336 18394 15369
rect 18235 15261 18267 15336
rect 18351 15261 18394 15336
rect 18235 15236 18394 15261
rect 23409 15324 23633 15368
rect 23409 15258 23462 15324
rect 23577 15258 23633 15324
rect 23409 15233 23633 15258
rect 27832 15334 28056 15371
rect 27832 15263 27888 15334
rect 28000 15263 28056 15334
rect 27832 15235 28056 15263
rect 32988 15339 33204 15360
rect 32988 15269 33040 15339
rect 33152 15269 33204 15339
rect 32988 15252 33204 15269
rect 35755 15333 35920 15357
rect 35755 15274 35784 15333
rect 35896 15274 35920 15333
rect 35755 15253 35920 15274
rect 45014 15136 46079 15485
rect 210 14825 296 14833
rect -1736 14821 296 14825
rect -1736 14765 224 14821
rect 280 14765 296 14821
rect -1736 14754 296 14765
rect -10148 12814 -2190 12867
rect -10148 12695 -2728 12814
rect -2419 12695 -2190 12814
rect -10148 12669 -2190 12695
rect -10148 7222 -7674 12669
rect -1736 9284 -1399 14754
rect 210 14750 296 14754
rect 2128 14495 2352 14515
rect 2128 14425 2184 14495
rect 2296 14425 2352 14495
rect 2128 14395 2352 14425
rect 6832 14489 7056 14515
rect 6832 14420 6888 14489
rect 7001 14420 7056 14489
rect 6832 14395 7056 14420
rect 11704 14494 11929 14515
rect 11704 14418 11760 14494
rect 11873 14418 11929 14494
rect 11704 14395 11929 14418
rect 16555 14478 16714 14499
rect 16555 14417 16592 14478
rect 16671 14417 16714 14478
rect 16555 14401 16714 14417
rect 21358 14481 21529 14504
rect 21358 14410 21397 14481
rect 21484 14410 21529 14481
rect 21358 14400 21529 14410
rect 26228 14483 26402 14503
rect 26228 14414 26265 14483
rect 26371 14414 26402 14483
rect 26228 14399 26402 14414
rect 31024 14479 31249 14498
rect 31024 14423 31080 14479
rect 31192 14423 31249 14479
rect 31024 14406 31249 14423
rect 37105 14489 37272 14508
rect 37105 14425 37150 14489
rect 37224 14425 37272 14489
rect 37105 14405 37272 14425
rect 2128 13383 2352 13403
rect 2128 13310 2184 13383
rect 2296 13310 2352 13383
rect 2128 13283 2352 13310
rect 6832 13374 7056 13403
rect 6832 13305 6885 13374
rect 7001 13305 7056 13374
rect 6832 13283 7056 13305
rect 11704 13384 11929 13402
rect 11704 13308 11760 13384
rect 11873 13308 11929 13384
rect 11704 13283 11929 13308
rect 16547 13372 16706 13392
rect 16547 13308 16594 13372
rect 16668 13308 16706 13372
rect 16547 13294 16706 13308
rect 21375 13376 21526 13393
rect 21375 13305 21406 13376
rect 21493 13305 21526 13376
rect 21375 13288 21526 13305
rect 26228 13380 26410 13396
rect 26228 13311 26267 13380
rect 26373 13311 26410 13380
rect 26228 13292 26410 13311
rect 31024 13370 31249 13390
rect 31024 13310 31080 13370
rect 31192 13310 31249 13370
rect 31024 13298 31249 13310
rect 37107 13376 37274 13394
rect 37107 13308 37148 13376
rect 37226 13308 37274 13376
rect 37107 13291 37274 13308
rect 48434 12843 50908 18233
rect -360 12825 50908 12843
rect -360 12824 37114 12825
rect -360 12822 6832 12824
rect -360 12708 -284 12822
rect -105 12809 6832 12822
rect -105 12708 2149 12809
rect -360 12689 2149 12708
rect 2320 12704 6832 12809
rect 7003 12819 37114 12824
rect 7003 12809 21367 12819
rect 7003 12805 16544 12809
rect 7003 12704 11721 12805
rect 2320 12689 11721 12704
rect -360 12685 11721 12689
rect 11892 12689 16544 12805
rect 16715 12699 21367 12809
rect 21538 12699 26218 12819
rect 26389 12814 37114 12819
rect 26389 12699 31032 12814
rect 16715 12694 31032 12699
rect 31203 12705 37114 12814
rect 37285 12705 50908 12825
rect 31203 12694 50908 12705
rect 16715 12689 50908 12694
rect 11892 12685 50908 12689
rect -360 12675 50908 12685
rect 45322 12671 50908 12675
rect 3807 12535 4033 12574
rect 363 12463 532 12498
rect 363 12402 396 12463
rect 501 12402 532 12463
rect 3807 12464 3864 12535
rect 3977 12464 4033 12535
rect 3807 12432 4033 12464
rect 8624 12549 8849 12574
rect 8624 12455 8681 12549
rect 8793 12455 8849 12549
rect 8624 12429 8849 12455
rect 13830 12535 14058 12579
rect 13830 12460 13885 12535
rect 14006 12460 14058 12535
rect 13830 12432 14058 12460
rect 18216 12530 18394 12566
rect 18216 12455 18268 12530
rect 18352 12455 18394 12530
rect 18216 12431 18394 12455
rect 23408 12526 23633 12555
rect 23408 12460 23462 12526
rect 23577 12460 23633 12526
rect 23408 12432 23633 12460
rect 27833 12527 28055 12559
rect 27833 12456 27889 12527
rect 28001 12456 28055 12527
rect 27833 12431 28055 12456
rect 33004 12535 33183 12558
rect 33004 12465 33040 12535
rect 33152 12465 33183 12535
rect 33004 12445 33183 12465
rect 35750 12524 35932 12542
rect 35750 12465 35784 12524
rect 35896 12465 35932 12524
rect 35750 12442 35932 12465
rect 363 12379 532 12402
rect 2128 11700 2352 11715
rect 2128 11616 2184 11700
rect 2296 11616 2352 11700
rect 2128 11595 2352 11616
rect 6832 11684 7056 11714
rect 6832 11615 6886 11684
rect 7002 11615 7056 11684
rect 6832 11594 7056 11615
rect 11704 11686 11929 11714
rect 11704 11611 11760 11686
rect 11872 11611 11929 11686
rect 11704 11595 11929 11611
rect 16567 11681 16716 11697
rect 16567 11617 16601 11681
rect 16675 11617 16716 11681
rect 16567 11603 16716 11617
rect 21365 11686 21516 11704
rect 21365 11610 21397 11686
rect 21483 11610 21516 11686
rect 21365 11599 21516 11610
rect 26230 11687 26412 11703
rect 26230 11611 26278 11687
rect 26367 11611 26412 11687
rect 26230 11599 26412 11611
rect 31024 11685 31248 11698
rect 31024 11625 31080 11685
rect 31192 11625 31248 11685
rect 31024 11610 31248 11625
rect 37094 11686 37270 11704
rect 37094 11618 37146 11686
rect 37224 11618 37270 11686
rect 37094 11603 37270 11618
rect 2128 10581 2352 10603
rect 2128 10503 2184 10581
rect 2296 10503 2352 10581
rect 2128 10483 2352 10503
rect 6831 10576 7055 10602
rect 6831 10505 6887 10576
rect 7001 10505 7055 10576
rect 6831 10482 7055 10505
rect 11704 10583 11928 10603
rect 11704 10508 11760 10583
rect 11872 10508 11928 10583
rect 11704 10483 11928 10508
rect 16560 10574 16709 10592
rect 16560 10512 16593 10574
rect 16669 10512 16709 10574
rect 16560 10498 16709 10512
rect 21357 10576 21525 10591
rect 21357 10500 21402 10576
rect 21488 10500 21525 10576
rect 21357 10489 21525 10500
rect 26228 10582 26415 10596
rect 26228 10506 26277 10582
rect 26366 10506 26415 10582
rect 26228 10489 26415 10506
rect 31024 10574 31248 10590
rect 31024 10518 31080 10574
rect 31193 10518 31248 10574
rect 31024 10502 31248 10518
rect 37093 10579 37269 10594
rect 37093 10506 37137 10579
rect 37219 10506 37269 10579
rect 37093 10493 37269 10506
rect 44997 10022 46321 10580
rect -367 9995 46321 10022
rect -367 9989 18215 9995
rect -367 9984 3841 9989
rect -367 9885 365 9984
rect 520 9890 3841 9984
rect 3996 9986 18215 9989
rect 3996 9890 8638 9986
rect 520 9887 8638 9890
rect 8793 9981 18215 9986
rect 8793 9887 13860 9981
rect 520 9885 13860 9887
rect -367 9882 13860 9885
rect 14015 9896 18215 9981
rect 18370 9993 46321 9995
rect 18370 9896 23449 9993
rect 14015 9894 23449 9896
rect 23604 9992 46321 9993
rect 23604 9981 33030 9992
rect 23604 9894 27863 9981
rect 14015 9882 27863 9894
rect 28018 9893 33030 9981
rect 33185 9981 46321 9992
rect 33185 9893 35753 9981
rect 28018 9882 35753 9893
rect 35908 9882 46321 9981
rect -367 9854 46321 9882
rect 336 9719 503 9744
rect 336 9654 368 9719
rect 474 9654 503 9719
rect 336 9632 503 9654
rect 3808 9741 4034 9767
rect 3808 9670 3863 9741
rect 3976 9670 4034 9741
rect 3808 9632 4034 9670
rect 8622 9730 8847 9762
rect 8622 9647 8680 9730
rect 8794 9647 8847 9730
rect 8622 9617 8847 9647
rect 13830 9735 14058 9780
rect 13830 9663 13887 9735
rect 14004 9663 14058 9735
rect 13830 9633 14058 9663
rect 18213 9735 18391 9766
rect 18213 9655 18265 9735
rect 18353 9655 18391 9735
rect 18213 9631 18391 9655
rect 23407 9726 23632 9763
rect 23407 9663 23463 9726
rect 23578 9663 23632 9726
rect 23407 9640 23632 9663
rect 27833 9733 28055 9762
rect 27833 9663 27888 9733
rect 28000 9663 28055 9733
rect 27833 9634 28055 9663
rect 33003 9732 33182 9760
rect 33003 9666 33031 9732
rect 33143 9666 33182 9732
rect 33003 9647 33182 9666
rect 35745 9732 35927 9755
rect 35745 9674 35784 9732
rect 35896 9674 35927 9732
rect 35745 9655 35927 9674
rect 44997 9380 46321 9854
rect 334 9284 419 9288
rect -1736 9278 419 9284
rect -1736 9214 344 9278
rect 408 9214 419 9278
rect -1736 9209 419 9214
rect -10148 7193 -2234 7222
rect -10148 7062 -2647 7193
rect -2418 7062 -2234 7193
rect -10148 7024 -2234 7062
rect -10148 1626 -7674 7024
rect -1736 6631 -1399 9209
rect 334 9203 419 9209
rect 2128 8893 2352 8915
rect 2128 8813 2184 8893
rect 2296 8813 2352 8893
rect 2128 8795 2352 8813
rect 6833 8885 7057 8913
rect 6833 8814 6886 8885
rect 7000 8814 7057 8885
rect 6833 8795 7057 8814
rect 11704 8889 11928 8914
rect 11704 8811 11760 8889
rect 11872 8811 11928 8889
rect 11704 8794 11928 8811
rect 16551 8878 16727 8900
rect 16551 8816 16598 8878
rect 16674 8816 16727 8878
rect 16551 8802 16727 8816
rect 21357 8885 21525 8904
rect 21357 8811 21397 8885
rect 21484 8811 21525 8885
rect 21357 8802 21525 8811
rect 26223 8886 26410 8907
rect 26223 8811 26265 8886
rect 26364 8811 26410 8886
rect 26223 8800 26410 8811
rect 31033 8882 31231 8900
rect 31033 8826 31079 8882
rect 31192 8826 31231 8882
rect 31033 8807 31231 8826
rect 37092 8885 37270 8901
rect 37092 8812 37142 8885
rect 37224 8812 37270 8885
rect 37092 8802 37270 8812
rect 2128 7784 2352 7803
rect 2128 7714 2184 7784
rect 2296 7714 2352 7784
rect 2128 7683 2352 7714
rect 6832 7773 7056 7802
rect 6832 7708 6888 7773
rect 7000 7708 7056 7773
rect 6832 7684 7056 7708
rect 11704 7781 11928 7802
rect 11704 7703 11760 7781
rect 11872 7703 11928 7781
rect 11704 7683 11928 7703
rect 16540 7772 16716 7791
rect 16540 7706 16589 7772
rect 16670 7706 16716 7772
rect 16540 7693 16716 7706
rect 21363 7779 21532 7793
rect 21363 7705 21404 7779
rect 21491 7705 21532 7779
rect 21363 7689 21532 7705
rect 26231 7783 26414 7796
rect 26231 7708 26273 7783
rect 26372 7708 26414 7783
rect 26231 7693 26414 7708
rect 31031 7772 31229 7790
rect 31031 7716 31079 7772
rect 31192 7716 31229 7772
rect 31031 7697 31229 7716
rect 37097 7779 37275 7794
rect 37097 7711 37144 7779
rect 37228 7711 37275 7779
rect 37097 7695 37275 7711
rect -382 7215 45449 7217
rect 48434 7215 50908 12671
rect -382 7208 50908 7215
rect -382 7190 26227 7208
rect -382 7188 11721 7190
rect -382 7066 -295 7188
rect -129 7185 11721 7188
rect -129 7180 6869 7185
rect -129 7066 2159 7180
rect -382 7060 2159 7066
rect 2330 7065 6869 7180
rect 7040 7070 11721 7185
rect 11892 7185 26227 7190
rect 11892 7070 16530 7185
rect 7040 7065 16530 7070
rect 16701 7180 26227 7185
rect 16701 7065 21334 7180
rect 2330 7060 21334 7065
rect 21505 7088 26227 7180
rect 26398 7194 50908 7208
rect 26398 7190 37088 7194
rect 26398 7088 31032 7190
rect 21505 7070 31032 7088
rect 31203 7074 37088 7190
rect 37259 7074 50908 7194
rect 31203 7070 50908 7074
rect 21505 7060 50908 7070
rect -382 7049 50908 7060
rect 45259 7043 50908 7049
rect 3807 6935 4033 6967
rect 337 6874 561 6900
rect 337 6805 390 6874
rect 505 6805 561 6874
rect 3807 6854 3863 6935
rect 3977 6854 4033 6935
rect 3807 6832 4033 6854
rect 8623 6928 8848 6965
rect 8623 6849 8679 6928
rect 8791 6849 8848 6928
rect 8623 6824 8848 6849
rect 13832 6938 14058 6973
rect 13832 6866 13886 6938
rect 14003 6866 14058 6938
rect 13832 6838 14058 6866
rect 18225 6956 18392 6977
rect 18225 6876 18263 6956
rect 18351 6876 18392 6956
rect 18225 6855 18392 6876
rect 23406 6928 23634 6962
rect 23406 6865 23462 6928
rect 23577 6865 23634 6928
rect 23406 6834 23634 6865
rect 27831 6939 28053 6967
rect 27831 6869 27887 6939
rect 27999 6869 28053 6939
rect 27831 6832 28053 6869
rect 33009 6930 33190 6951
rect 33009 6864 33041 6930
rect 33153 6864 33190 6930
rect 33009 6842 33190 6864
rect 35737 6921 35937 6945
rect 35737 6863 35784 6921
rect 35896 6863 35937 6921
rect 35737 6839 35937 6863
rect 337 6779 561 6805
rect -1736 6559 621 6631
rect -1736 3684 -1399 6559
rect 549 6489 621 6559
rect 544 6479 628 6489
rect 544 6416 554 6479
rect 618 6416 628 6479
rect 544 6406 628 6416
rect 2128 6088 2352 6115
rect 2128 6012 2184 6088
rect 2296 6012 2352 6088
rect 2128 5995 2352 6012
rect 6832 6081 7056 6115
rect 6832 6016 6888 6081
rect 7000 6016 7056 6081
rect 6832 5995 7056 6016
rect 11703 6089 11927 6114
rect 11703 6016 11761 6089
rect 11874 6016 11927 6089
rect 11703 5995 11927 6016
rect 16558 6082 16730 6104
rect 16558 6016 16593 6082
rect 16674 6016 16730 6082
rect 16558 5998 16730 6016
rect 21359 6083 21528 6105
rect 21359 6011 21400 6083
rect 21485 6011 21528 6083
rect 21359 6001 21528 6011
rect 26232 6090 26415 6102
rect 26232 6010 26275 6090
rect 26367 6010 26415 6090
rect 26232 5999 26415 6010
rect 31049 6082 31220 6098
rect 31049 6026 31080 6082
rect 31193 6026 31220 6082
rect 31049 6009 31220 6026
rect 37090 6083 37270 6101
rect 37090 6015 37140 6083
rect 37224 6015 37270 6083
rect 37090 6002 37270 6015
rect 2128 4984 2353 5003
rect 2128 4910 2184 4984
rect 2296 4910 2353 4984
rect 2128 4883 2353 4910
rect 6832 4974 7056 5003
rect 6832 4903 6888 4974
rect 7001 4903 7056 4974
rect 6832 4883 7056 4903
rect 11704 4980 11929 5002
rect 11704 4907 11759 4980
rect 11872 4907 11929 4980
rect 11704 4883 11929 4907
rect 16545 4976 16717 4993
rect 16545 4906 16589 4976
rect 16672 4906 16717 4976
rect 16545 4887 16717 4906
rect 21375 4974 21532 4993
rect 21375 4902 21408 4974
rect 21493 4902 21532 4974
rect 21375 4887 21532 4902
rect 26242 4980 26415 4996
rect 26242 4900 26281 4980
rect 26373 4900 26415 4980
rect 31050 4977 31221 4990
rect 31050 4921 31080 4977
rect 31192 4921 31221 4977
rect 31050 4901 31221 4921
rect 37100 4976 37280 4992
rect 37100 4910 37140 4976
rect 37228 4910 37280 4976
rect 26242 4886 26415 4900
rect 37100 4893 37280 4910
rect 45047 4433 46330 5073
rect -338 4417 46330 4433
rect -338 4413 8638 4417
rect -338 4307 359 4413
rect 523 4376 8638 4413
rect 523 4307 3830 4376
rect -338 4270 3830 4307
rect 3994 4311 8638 4376
rect 8802 4403 46330 4417
rect 8802 4397 35760 4403
rect 8802 4392 18225 4397
rect 8802 4311 13830 4392
rect 3994 4286 13830 4311
rect 13994 4291 18225 4392
rect 18389 4291 23429 4397
rect 23593 4291 27849 4397
rect 28013 4392 35760 4397
rect 28013 4291 33020 4392
rect 13994 4286 33020 4291
rect 33184 4297 35760 4392
rect 35924 4297 46330 4403
rect 33184 4286 46330 4297
rect 3994 4270 46330 4286
rect -338 4265 46330 4270
rect 336 4141 561 4200
rect 336 4062 390 4141
rect 507 4062 561 4141
rect 336 4028 561 4062
rect 3808 4139 4032 4172
rect 3808 4058 3863 4139
rect 3977 4058 4032 4139
rect 3808 4031 4032 4058
rect 8624 4129 8849 4164
rect 8624 4052 8680 4129
rect 8793 4052 8849 4129
rect 8624 4025 8849 4052
rect 13831 4135 14057 4166
rect 13831 4060 13887 4135
rect 14000 4060 14057 4135
rect 13831 4033 14057 4060
rect 18222 4141 18389 4170
rect 18222 4066 18267 4141
rect 18360 4066 18389 4141
rect 18222 4048 18389 4066
rect 23407 4127 23635 4161
rect 23407 4056 23460 4127
rect 23576 4056 23635 4127
rect 23407 4033 23635 4056
rect 27834 4123 28056 4160
rect 27834 4050 27887 4123
rect 28001 4050 28056 4123
rect 27834 4025 28056 4050
rect 32997 4136 33178 4158
rect 32997 4072 33030 4136
rect 33139 4072 33178 4136
rect 32997 4049 33178 4072
rect 35742 4130 35942 4159
rect 35742 4074 35783 4130
rect 35896 4074 35942 4130
rect 35742 4053 35942 4074
rect 45047 3809 46330 4265
rect 318 3684 401 3687
rect -1736 3677 401 3684
rect -1736 3617 328 3677
rect 391 3617 401 3677
rect -1736 3614 401 3617
rect -1736 2800 -1399 3614
rect 318 3607 401 3614
rect 2128 3293 2352 3315
rect 2128 3214 2184 3293
rect 2296 3214 2352 3293
rect 2128 3195 2352 3214
rect 6832 3288 7056 3314
rect 6832 3217 6888 3288
rect 7001 3217 7056 3288
rect 6832 3194 7056 3217
rect 11701 3284 11926 3314
rect 11701 3209 11757 3284
rect 11875 3209 11926 3284
rect 11701 3195 11926 3209
rect 16560 3288 16719 3302
rect 16560 3218 16594 3288
rect 16677 3218 16719 3288
rect 16560 3202 16719 3218
rect 21371 3283 21528 3303
rect 21371 3212 21401 3283
rect 21486 3212 21528 3283
rect 21371 3197 21528 3212
rect 26229 3290 26402 3309
rect 26229 3210 26264 3290
rect 26360 3210 26402 3290
rect 26229 3199 26402 3210
rect 31051 3278 31233 3299
rect 31051 3222 31080 3278
rect 31192 3222 31233 3278
rect 31051 3204 31233 3222
rect 37093 3285 37278 3305
rect 37093 3219 37137 3285
rect 37225 3219 37278 3285
rect 37093 3206 37278 3219
rect 2128 2172 2352 2203
rect 2128 2104 2184 2172
rect 2296 2104 2352 2172
rect 2128 2083 2352 2104
rect 6832 2173 7056 2204
rect 6832 2104 6887 2173
rect 7001 2104 7056 2173
rect 6832 2084 7056 2104
rect 11702 2181 11929 2200
rect 11702 2106 11758 2181
rect 11876 2106 11929 2181
rect 11702 2085 11929 2106
rect 16553 2177 16712 2194
rect 16553 2104 16595 2177
rect 16675 2104 16712 2177
rect 16553 2094 16712 2104
rect 21376 2174 21524 2196
rect 21376 2103 21403 2174
rect 21488 2103 21524 2174
rect 21376 2084 21524 2103
rect 26227 2179 26412 2195
rect 26227 2099 26276 2179
rect 26372 2099 26412 2179
rect 31046 2178 31228 2194
rect 31046 2117 31079 2178
rect 31193 2117 31228 2178
rect 31046 2099 31228 2117
rect 26227 2088 26412 2099
rect -10148 1620 687 1626
rect 21225 1620 22014 1621
rect 30989 1620 31336 1621
rect 37039 1620 37388 1759
rect -10148 1616 45603 1620
rect 48434 1616 50908 7043
rect -10148 1601 50908 1616
rect -10148 1481 2140 1601
rect 2311 1597 50908 1601
rect 2311 1596 37103 1597
rect 2311 1591 16552 1596
rect 2311 1587 11691 1591
rect 2311 1481 6848 1587
rect -10148 1467 6848 1481
rect 7019 1471 11691 1587
rect 11862 1476 16552 1591
rect 16723 1595 37103 1596
rect 16723 1591 31033 1595
rect 16723 1576 26229 1591
rect 16723 1486 21377 1576
rect 21510 1486 26229 1576
rect 16723 1476 26229 1486
rect 11862 1471 26229 1476
rect 26400 1475 31033 1591
rect 31204 1477 37103 1595
rect 37274 1477 50908 1597
rect 31204 1475 50908 1477
rect 26400 1471 50908 1475
rect 7019 1467 50908 1471
rect -10148 1452 50908 1467
rect -10148 1451 687 1452
rect -10148 -4926 -7674 1451
rect 2062 520 2406 1452
rect 3808 1332 4032 1378
rect 3808 1265 3864 1332
rect 3976 1265 4032 1332
rect 3808 1232 4032 1265
rect 6783 603 7127 1452
rect 8625 1334 8849 1364
rect 8625 1257 8679 1334
rect 8792 1257 8849 1334
rect 8625 1231 8849 1257
rect 2061 489 2410 520
rect 2061 416 2184 489
rect 2296 416 2410 489
rect 2061 -4926 2410 416
rect 6778 487 7127 603
rect 11646 578 11990 1452
rect 13834 1328 14055 1363
rect 13834 1255 13872 1328
rect 14002 1255 14055 1328
rect 13834 1219 14055 1255
rect 6778 418 6887 487
rect 7001 418 7127 487
rect 6778 -4926 7127 418
rect 11645 487 11994 578
rect 16467 566 16811 1452
rect 21225 1451 22014 1452
rect 18198 1335 18424 1361
rect 18198 1260 18262 1335
rect 18355 1260 18424 1335
rect 18198 1233 18424 1260
rect 21276 689 21624 1451
rect 23409 1342 23632 1368
rect 23409 1271 23462 1342
rect 23578 1271 23632 1342
rect 23409 1233 23632 1271
rect 26160 720 26506 1452
rect 27832 1330 28059 1357
rect 27832 1257 27887 1330
rect 28001 1257 28059 1330
rect 27832 1233 28059 1257
rect 30989 775 31336 1452
rect 33008 1329 33186 1356
rect 33008 1265 33043 1329
rect 33152 1265 33186 1329
rect 33008 1241 33186 1265
rect 11645 410 11760 487
rect 11872 410 11994 487
rect 11645 -4926 11994 410
rect 16463 485 16812 566
rect 16463 412 16588 485
rect 16668 412 16812 485
rect 16463 -4926 16812 412
rect 21276 480 21625 689
rect 21276 408 21402 480
rect 21481 408 21625 480
rect 21276 -4926 21625 408
rect 26159 483 26508 720
rect 26159 406 26275 483
rect 26363 406 26508 483
rect 26159 -4926 26508 406
rect 30986 521 31336 775
rect 30986 482 31335 521
rect 30986 421 31079 482
rect 31193 421 31335 482
rect 30986 -4926 31335 421
rect 37039 -4926 37388 1452
rect 45385 1444 50908 1452
rect 48434 -4926 50908 1444
rect -10148 -7521 50920 -4926
rect -10147 -7526 50920 -7521
<< via3 >>
rect 2120 27854 2373 28125
rect 6889 27707 7064 27952
rect 11691 28067 11959 28436
rect 16525 28225 16765 28508
rect 21331 28222 21592 28583
rect 26205 27940 26457 28269
rect 31016 28204 31278 28484
rect 35784 27796 35874 27869
rect 40384 29049 40502 29131
rect 37124 27023 37213 27079
rect 35801 26846 35890 26918
rect 37123 26063 37244 26128
rect 35794 25881 35883 25953
rect 37126 25104 37244 25163
rect 35800 24915 35893 24993
rect 391 22657 504 22733
rect 8680 23169 8793 23243
rect 13888 23184 13944 23240
rect 18283 23184 18339 23240
rect 23493 23184 23549 23240
rect 27862 23179 28000 23251
rect 37119 24130 37237 24189
rect 3881 22614 3971 22672
rect 11761 22389 11874 22465
rect 16605 22400 16661 22456
rect 21421 22400 21477 22456
rect 26292 22400 26348 22456
rect 31111 22400 31167 22456
rect 2184 21703 2296 21777
rect 6887 21698 7001 21776
rect 11760 21700 11873 21782
rect 16593 21710 16683 21769
rect 21412 21709 21490 21773
rect 26264 21706 26375 21776
rect 31080 21714 31193 21771
rect 37146 21707 37224 21773
rect -3218 18260 -3023 18392
rect 402 21105 487 21181
rect 3887 21103 3972 21179
rect 8706 21103 8791 21179
rect 13893 21097 13978 21173
rect 18269 21103 18354 21179
rect 23473 21097 23558 21173
rect 27903 21109 27988 21185
rect 33024 21097 33109 21173
rect 35797 21099 35882 21175
rect 392 20849 505 20925
rect 3864 20871 3976 20940
rect 8678 20855 8793 20940
rect 13889 20866 14003 20934
rect 18268 20864 18348 20943
rect 23462 20862 23576 20944
rect 27887 20864 28000 20937
rect 33039 20874 33155 20938
rect 35784 20869 35896 20928
rect 2184 20019 2296 20085
rect 6888 20014 7000 20091
rect 11760 20016 11872 20098
rect 16583 20022 16673 20081
rect 21409 20021 21486 20085
rect 26277 20017 26366 20089
rect 31079 20020 31192 20077
rect 37145 20023 37223 20089
rect 2184 18907 2296 18973
rect 6888 18901 7000 18976
rect 11760 18904 11872 18986
rect 16593 18910 16665 18969
rect 21404 18914 21481 18978
rect 26281 18903 26370 18975
rect 31080 18911 31192 18969
rect 37151 18909 37227 18978
rect -217 18265 -32 18368
rect 2155 18258 2326 18368
rect 6871 18264 7042 18374
rect 11718 18270 11889 18380
rect 16548 18258 16719 18368
rect 21374 18262 21545 18382
rect 26231 18254 26402 18374
rect 31048 18258 31219 18378
rect 37093 18254 37264 18374
rect 392 18005 505 18072
rect 3863 18059 3977 18136
rect 8680 18055 8792 18139
rect 13888 18070 14002 18138
rect 18269 18065 18349 18144
rect 23464 18068 23575 18143
rect 27889 18066 28002 18139
rect 33038 18053 33154 18117
rect 35784 18068 35896 18127
rect 2184 17214 2296 17300
rect 6888 17221 7000 17291
rect 11761 17212 11872 17282
rect 16599 17219 16671 17278
rect 21407 17212 21487 17285
rect 26270 17214 26369 17285
rect 31080 17221 31192 17279
rect 37143 17220 37219 17289
rect 2184 16117 2296 16181
rect 6887 16104 7000 16173
rect 11762 16110 11873 16180
rect 16588 16114 16667 16175
rect 21411 16108 21491 16181
rect 26271 16105 26370 16176
rect 31080 16115 31192 16171
rect 37144 16111 37218 16175
rect 439 15539 503 15603
rect 3877 15529 3941 15593
rect 8694 15529 8758 15593
rect 13902 15529 13966 15593
rect 18260 15534 18324 15598
rect 23473 15534 23537 15598
rect 27903 15536 27967 15600
rect 33057 15541 33121 15605
rect 35802 15544 35866 15608
rect 378 15254 513 15321
rect 3863 15255 3977 15332
rect 8679 15249 8791 15343
rect 13887 15263 14008 15338
rect 18267 15261 18351 15336
rect 23462 15258 23577 15324
rect 33040 15269 33152 15339
rect 35784 15274 35896 15333
rect -2728 12695 -2419 12814
rect 2184 14425 2296 14495
rect 6888 14420 7001 14489
rect 11760 14418 11873 14494
rect 16592 14417 16671 14478
rect 21397 14410 21484 14481
rect 26265 14414 26371 14483
rect 31080 14423 31192 14479
rect 37150 14425 37224 14489
rect 2184 13310 2296 13383
rect 6885 13305 7001 13374
rect 11760 13308 11873 13384
rect 16594 13308 16668 13372
rect 21406 13305 21493 13376
rect 26267 13311 26373 13380
rect 31080 13310 31192 13370
rect 37148 13308 37226 13376
rect -284 12708 -105 12822
rect 2149 12689 2320 12809
rect 6832 12704 7003 12824
rect 11721 12685 11892 12805
rect 16544 12689 16715 12809
rect 21367 12699 21538 12819
rect 26218 12699 26389 12819
rect 31032 12694 31203 12814
rect 37114 12705 37285 12825
rect 396 12402 501 12463
rect 3864 12464 3977 12535
rect 8681 12455 8793 12549
rect 13885 12460 14006 12535
rect 18268 12455 18352 12530
rect 23462 12460 23577 12526
rect 27889 12456 28001 12527
rect 33040 12465 33152 12535
rect 35784 12465 35896 12524
rect 2184 11616 2296 11700
rect 6886 11615 7002 11684
rect 11760 11611 11872 11686
rect 16601 11617 16675 11681
rect 21397 11610 21483 11686
rect 26278 11611 26367 11687
rect 31080 11625 31192 11685
rect 37146 11618 37224 11686
rect 2184 10503 2296 10581
rect 6887 10505 7001 10576
rect 11760 10508 11872 10583
rect 16593 10512 16669 10574
rect 21402 10500 21488 10576
rect 26277 10506 26366 10582
rect 31080 10518 31193 10574
rect 37137 10506 37219 10579
rect 365 9885 520 9984
rect 3841 9890 3996 9989
rect 8638 9887 8793 9986
rect 13860 9882 14015 9981
rect 18215 9896 18370 9995
rect 23449 9894 23604 9993
rect 27863 9882 28018 9981
rect 33030 9893 33185 9992
rect 35753 9882 35908 9981
rect 368 9654 474 9719
rect 3863 9670 3976 9741
rect 8680 9647 8794 9730
rect 13887 9663 14004 9735
rect 18265 9655 18353 9735
rect 23463 9663 23578 9726
rect 27888 9663 28000 9733
rect 33031 9666 33143 9732
rect 35784 9674 35896 9732
rect -2647 7062 -2418 7193
rect 2184 8813 2296 8893
rect 6886 8814 7000 8885
rect 11760 8811 11872 8889
rect 16598 8816 16674 8878
rect 21397 8811 21484 8885
rect 26265 8811 26364 8886
rect 31079 8826 31192 8882
rect 37142 8812 37224 8885
rect 2184 7714 2296 7784
rect 6888 7708 7000 7773
rect 11760 7703 11872 7781
rect 16589 7706 16670 7772
rect 21404 7705 21491 7779
rect 26273 7708 26372 7783
rect 31079 7716 31192 7772
rect 37144 7711 37228 7779
rect -295 7066 -129 7188
rect 2159 7060 2330 7180
rect 6869 7065 7040 7185
rect 11721 7070 11892 7190
rect 16530 7065 16701 7185
rect 21334 7060 21505 7180
rect 26227 7088 26398 7208
rect 31032 7070 31203 7190
rect 37088 7074 37259 7194
rect 390 6805 505 6874
rect 3863 6854 3977 6935
rect 8679 6849 8791 6928
rect 13886 6866 14003 6938
rect 18263 6876 18351 6956
rect 23462 6865 23577 6928
rect 33041 6864 33153 6930
rect 35784 6863 35896 6921
rect 2184 6012 2296 6088
rect 6888 6016 7000 6081
rect 11761 6016 11874 6089
rect 16593 6016 16674 6082
rect 21400 6011 21485 6083
rect 26275 6010 26367 6090
rect 31080 6026 31193 6082
rect 37140 6015 37224 6083
rect 2184 4910 2296 4984
rect 6888 4903 7001 4974
rect 11759 4907 11872 4980
rect 16589 4906 16672 4976
rect 21408 4902 21493 4974
rect 26281 4900 26373 4980
rect 31080 4921 31192 4977
rect 37140 4910 37228 4976
rect 359 4307 523 4413
rect 3830 4270 3994 4376
rect 8638 4311 8802 4417
rect 13830 4286 13994 4392
rect 18225 4291 18389 4397
rect 23429 4291 23593 4397
rect 27849 4291 28013 4397
rect 33020 4286 33184 4392
rect 35760 4297 35924 4403
rect 390 4062 507 4141
rect 3863 4058 3977 4139
rect 8680 4052 8793 4129
rect 13887 4060 14000 4135
rect 18267 4066 18360 4141
rect 23460 4056 23576 4127
rect 27887 4050 28001 4123
rect 33030 4072 33139 4136
rect 35783 4074 35896 4130
rect 2184 3214 2296 3293
rect 6888 3217 7001 3288
rect 11757 3209 11875 3284
rect 16594 3218 16677 3288
rect 21401 3212 21486 3283
rect 26264 3210 26360 3290
rect 31080 3222 31192 3278
rect 37137 3219 37225 3285
rect 2184 2104 2296 2172
rect 6887 2104 7001 2173
rect 11758 2106 11876 2181
rect 16595 2104 16675 2177
rect 21403 2103 21488 2174
rect 26276 2099 26372 2179
rect 31079 2117 31193 2178
rect 2140 1481 2311 1601
rect 6848 1467 7019 1587
rect 11691 1471 11862 1591
rect 16552 1476 16723 1596
rect 21377 1486 21510 1576
rect 26229 1471 26400 1591
rect 31033 1475 31204 1595
rect 37103 1477 37274 1597
rect 3864 1265 3976 1332
rect 8679 1257 8792 1334
rect 2184 416 2296 489
rect 13872 1255 14002 1328
rect 6887 418 7001 487
rect 18262 1260 18355 1335
rect 23462 1271 23578 1342
rect 27887 1257 28001 1330
rect 33043 1265 33152 1329
rect 11760 410 11872 487
rect 16588 412 16668 485
rect 21402 408 21481 480
rect 26275 406 26363 483
rect 31079 421 31193 482
<< metal4 >>
rect 44398 32676 46994 32701
rect -6208 30269 46994 32676
rect -6233 30206 46994 30269
rect -6233 30202 47058 30206
rect -6233 21224 -3581 30202
rect 293 27719 649 30202
rect 280 27310 649 27719
rect 2070 28125 2417 28254
rect 2070 27854 2120 28125
rect 2373 27854 2417 28125
rect 280 22733 616 27310
rect 280 22657 391 22733
rect 504 22657 616 22733
rect 280 22260 616 22657
rect 311 22120 616 22260
rect 280 21516 616 22120
rect 2070 21938 2417 27854
rect 3727 27719 4083 30202
rect 6775 27952 7122 28174
rect 3727 27175 4088 27719
rect 3752 22672 4088 27175
rect 3752 22614 3881 22672
rect 3971 22614 4088 22672
rect 281 21366 616 21516
rect 280 21224 616 21366
rect -6233 21181 616 21224
rect -6233 21105 402 21181
rect 487 21105 616 21181
rect -6233 21047 616 21105
rect -6233 15695 -3581 21047
rect 280 20925 616 21047
rect 280 20849 392 20925
rect 505 20849 616 20925
rect -3290 18392 85 18408
rect -3290 18260 -3218 18392
rect -3023 18368 85 18392
rect -3023 18265 -217 18368
rect -32 18265 85 18368
rect -3023 18260 85 18265
rect -3290 18237 85 18260
rect 280 18072 616 20849
rect 280 18005 392 18072
rect 505 18005 616 18072
rect 280 15695 616 18005
rect -6233 15603 616 15695
rect -6233 15539 439 15603
rect 503 15539 616 15603
rect -6233 15428 616 15539
rect -6233 10087 -3581 15428
rect 280 15321 616 15428
rect 280 15254 378 15321
rect 513 15254 616 15321
rect -2850 12822 -44 12847
rect -2850 12814 -284 12822
rect -2850 12695 -2728 12814
rect -2419 12708 -284 12814
rect -105 12708 -44 12822
rect -2419 12695 -44 12708
rect -2850 12676 -44 12695
rect 280 12463 616 15254
rect 280 12402 396 12463
rect 501 12402 616 12463
rect 280 10087 616 12402
rect -6233 9984 616 10087
rect -6233 9885 365 9984
rect 520 9885 616 9984
rect -6233 9820 616 9885
rect -6233 4480 -3581 9820
rect 280 9719 616 9820
rect 280 9654 368 9719
rect 474 9654 616 9719
rect -2899 7193 14 7217
rect -2899 7062 -2647 7193
rect -2418 7188 14 7193
rect -2418 7066 -295 7188
rect -129 7066 14 7188
rect -2418 7062 14 7066
rect -2899 7046 14 7062
rect 280 6874 616 9654
rect 280 6805 390 6874
rect 505 6805 616 6874
rect 280 4480 616 6805
rect -6233 4413 616 4480
rect -6233 4307 359 4413
rect 523 4307 616 4413
rect -6233 4213 616 4307
rect -6233 -1009 -3581 4213
rect 280 4141 616 4213
rect 280 4062 390 4141
rect 507 4062 616 4141
rect 280 699 616 4062
rect 2072 21777 2408 21938
rect 2072 21703 2184 21777
rect 2296 21703 2408 21777
rect 2072 20085 2408 21703
rect 2072 20019 2184 20085
rect 2296 20019 2408 20085
rect 2072 18973 2408 20019
rect 2072 18907 2184 18973
rect 2296 18907 2408 18973
rect 2072 18368 2408 18907
rect 2072 18258 2155 18368
rect 2326 18258 2408 18368
rect 2072 17300 2408 18258
rect 2072 17214 2184 17300
rect 2296 17214 2408 17300
rect 2072 16181 2408 17214
rect 2072 16117 2184 16181
rect 2296 16117 2408 16181
rect 2072 14495 2408 16117
rect 2072 14425 2184 14495
rect 2296 14425 2408 14495
rect 2072 13383 2408 14425
rect 2072 13310 2184 13383
rect 2296 13310 2408 13383
rect 2072 12809 2408 13310
rect 2072 12689 2149 12809
rect 2320 12689 2408 12809
rect 2072 11700 2408 12689
rect 2072 11616 2184 11700
rect 2296 11616 2408 11700
rect 2072 10581 2408 11616
rect 2072 10503 2184 10581
rect 2296 10503 2408 10581
rect 2072 8893 2408 10503
rect 2072 8813 2184 8893
rect 2296 8813 2408 8893
rect 2072 7784 2408 8813
rect 2072 7714 2184 7784
rect 2296 7714 2408 7784
rect 2072 7180 2408 7714
rect 2072 7060 2159 7180
rect 2330 7060 2408 7180
rect 2072 6088 2408 7060
rect 2072 6012 2184 6088
rect 2296 6012 2408 6088
rect 2072 4984 2408 6012
rect 2072 4910 2184 4984
rect 2296 4910 2408 4984
rect 2072 3293 2408 4910
rect 2072 3214 2184 3293
rect 2296 3214 2408 3293
rect 2072 2172 2408 3214
rect 2072 2104 2184 2172
rect 2296 2104 2408 2172
rect 2072 1601 2408 2104
rect 2072 1481 2140 1601
rect 2311 1481 2408 1601
rect 275 -1002 617 699
rect 2072 489 2408 1481
rect 2072 416 2184 489
rect 2296 416 2408 489
rect 2072 305 2408 416
rect 2069 168 2408 305
rect 3752 21179 4088 22614
rect 6775 27707 6889 27952
rect 7064 27707 7122 27952
rect 6775 21858 7122 27707
rect 8557 27238 8913 30202
rect 11647 28436 11994 29111
rect 11647 28067 11691 28436
rect 11959 28067 11994 28436
rect 8568 23243 8904 27238
rect 8568 23169 8680 23243
rect 8793 23169 8904 23243
rect 3752 21103 3887 21179
rect 3972 21103 4088 21179
rect 3752 20940 4088 21103
rect 3752 20871 3864 20940
rect 3976 20871 4088 20940
rect 3752 18136 4088 20871
rect 3752 18059 3863 18136
rect 3977 18059 4088 18136
rect 3752 15593 4088 18059
rect 3752 15529 3877 15593
rect 3941 15529 4088 15593
rect 3752 15332 4088 15529
rect 3752 15255 3863 15332
rect 3977 15255 4088 15332
rect 3752 12535 4088 15255
rect 3752 12464 3864 12535
rect 3977 12464 4088 12535
rect 3752 9989 4088 12464
rect 3752 9890 3841 9989
rect 3996 9890 4088 9989
rect 3752 9741 4088 9890
rect 3752 9670 3863 9741
rect 3976 9670 4088 9741
rect 3752 6935 4088 9670
rect 3752 6854 3863 6935
rect 3977 6854 4088 6935
rect 3752 4376 4088 6854
rect 3752 4270 3830 4376
rect 3994 4270 4088 4376
rect 3752 4139 4088 4270
rect 3752 4058 3863 4139
rect 3977 4058 4088 4139
rect 3752 1332 4088 4058
rect 3752 1265 3864 1332
rect 3976 1265 4088 1332
rect 3752 230 4088 1265
rect 3751 168 4088 230
rect 6776 21776 7112 21858
rect 6776 21698 6887 21776
rect 7001 21698 7112 21776
rect 6776 20091 7112 21698
rect 6776 20014 6888 20091
rect 7000 20014 7112 20091
rect 6776 18976 7112 20014
rect 6776 18901 6888 18976
rect 7000 18901 7112 18976
rect 6776 18374 7112 18901
rect 6776 18264 6871 18374
rect 7042 18264 7112 18374
rect 6776 17291 7112 18264
rect 6776 17221 6888 17291
rect 7000 17221 7112 17291
rect 6776 16173 7112 17221
rect 6776 16104 6887 16173
rect 7000 16104 7112 16173
rect 6776 14489 7112 16104
rect 6776 14420 6888 14489
rect 7001 14420 7112 14489
rect 6776 13374 7112 14420
rect 6776 13305 6885 13374
rect 7001 13305 7112 13374
rect 6776 12824 7112 13305
rect 6776 12704 6832 12824
rect 7003 12704 7112 12824
rect 6776 11684 7112 12704
rect 6776 11615 6886 11684
rect 7002 11615 7112 11684
rect 6776 10576 7112 11615
rect 6776 10505 6887 10576
rect 7001 10505 7112 10576
rect 6776 8885 7112 10505
rect 6776 8814 6886 8885
rect 7000 8814 7112 8885
rect 6776 7773 7112 8814
rect 6776 7708 6888 7773
rect 7000 7708 7112 7773
rect 6776 7185 7112 7708
rect 6776 7065 6869 7185
rect 7040 7065 7112 7185
rect 6776 6081 7112 7065
rect 6776 6016 6888 6081
rect 7000 6016 7112 6081
rect 6776 4974 7112 6016
rect 6776 4903 6888 4974
rect 7001 4903 7112 4974
rect 6776 3288 7112 4903
rect 6776 3217 6888 3288
rect 7001 3217 7112 3288
rect 6776 2173 7112 3217
rect 6776 2104 6887 2173
rect 7001 2104 7112 2173
rect 6776 1587 7112 2104
rect 6776 1467 6848 1587
rect 7019 1467 7112 1587
rect 6776 487 7112 1467
rect 6776 418 6887 487
rect 7001 418 7112 487
rect 2069 -252 2406 168
rect 2069 -711 2404 -252
rect 3751 -1002 4085 168
rect 6776 0 7112 418
rect 8568 21179 8904 23169
rect 11647 22795 11994 28067
rect 13775 27382 14131 30202
rect 16460 28508 16807 28892
rect 16460 28225 16525 28508
rect 16765 28225 16807 28508
rect 13776 23240 14112 27382
rect 13776 23184 13888 23240
rect 13944 23184 14112 23240
rect 8568 21103 8706 21179
rect 8791 21103 8904 21179
rect 8568 20940 8904 21103
rect 8568 20855 8678 20940
rect 8793 20855 8904 20940
rect 8568 18139 8904 20855
rect 8568 18055 8680 18139
rect 8792 18055 8904 18139
rect 8568 15593 8904 18055
rect 8568 15529 8694 15593
rect 8758 15529 8904 15593
rect 8568 15343 8904 15529
rect 8568 15249 8679 15343
rect 8791 15249 8904 15343
rect 8568 12549 8904 15249
rect 8568 12455 8681 12549
rect 8793 12455 8904 12549
rect 8568 9986 8904 12455
rect 8568 9887 8638 9986
rect 8793 9887 8904 9986
rect 8568 9730 8904 9887
rect 8568 9647 8680 9730
rect 8794 9647 8904 9730
rect 8568 6928 8904 9647
rect 8568 6849 8679 6928
rect 8791 6849 8904 6928
rect 8568 4417 8904 6849
rect 8568 4311 8638 4417
rect 8802 4311 8904 4417
rect 8568 4129 8904 4311
rect 8568 4052 8680 4129
rect 8793 4052 8904 4129
rect 8568 1334 8904 4052
rect 8568 1257 8679 1334
rect 8792 1257 8904 1334
rect 8568 56 8904 1257
rect 11648 22465 11984 22795
rect 11648 22389 11761 22465
rect 11874 22389 11984 22465
rect 11648 21782 11984 22389
rect 11648 21700 11760 21782
rect 11873 21700 11984 21782
rect 11648 20098 11984 21700
rect 11648 20016 11760 20098
rect 11872 20016 11984 20098
rect 11648 18986 11984 20016
rect 11648 18904 11760 18986
rect 11872 18904 11984 18986
rect 11648 18380 11984 18904
rect 11648 18270 11718 18380
rect 11889 18270 11984 18380
rect 11648 17282 11984 18270
rect 11648 17212 11761 17282
rect 11872 17212 11984 17282
rect 11648 16180 11984 17212
rect 11648 16110 11762 16180
rect 11873 16110 11984 16180
rect 11648 14494 11984 16110
rect 11648 14418 11760 14494
rect 11873 14418 11984 14494
rect 11648 13384 11984 14418
rect 11648 13308 11760 13384
rect 11873 13308 11984 13384
rect 11648 12805 11984 13308
rect 11648 12685 11721 12805
rect 11892 12685 11984 12805
rect 11648 11686 11984 12685
rect 11648 11611 11760 11686
rect 11872 11611 11984 11686
rect 11648 10583 11984 11611
rect 11648 10508 11760 10583
rect 11872 10508 11984 10583
rect 11648 8889 11984 10508
rect 11648 8811 11760 8889
rect 11872 8811 11984 8889
rect 11648 7781 11984 8811
rect 11648 7703 11760 7781
rect 11872 7703 11984 7781
rect 11648 7190 11984 7703
rect 11648 7070 11721 7190
rect 11892 7070 11984 7190
rect 11648 6089 11984 7070
rect 11648 6016 11761 6089
rect 11874 6016 11984 6089
rect 11648 4980 11984 6016
rect 11648 4907 11759 4980
rect 11872 4907 11984 4980
rect 11648 3284 11984 4907
rect 11648 3209 11757 3284
rect 11875 3209 11984 3284
rect 11648 2181 11984 3209
rect 13776 21173 14112 23184
rect 16460 22576 16807 28225
rect 18137 27319 18493 30202
rect 21284 28583 21631 28918
rect 21284 28222 21331 28583
rect 21592 28222 21631 28583
rect 18144 24528 18480 27319
rect 18144 23240 18481 24528
rect 18144 23184 18283 23240
rect 18339 23184 18481 23240
rect 13776 21097 13893 21173
rect 13978 21097 14112 21173
rect 13776 20934 14112 21097
rect 13776 20866 13889 20934
rect 14003 20866 14112 20934
rect 13776 18138 14112 20866
rect 13776 18070 13888 18138
rect 14002 18070 14112 18138
rect 13776 15593 14112 18070
rect 13776 15529 13902 15593
rect 13966 15529 14112 15593
rect 13776 15338 14112 15529
rect 13776 15263 13887 15338
rect 14008 15263 14112 15338
rect 13776 12535 14112 15263
rect 13776 12460 13885 12535
rect 14006 12460 14112 12535
rect 13776 9981 14112 12460
rect 13776 9882 13860 9981
rect 14015 9882 14112 9981
rect 13776 9735 14112 9882
rect 13776 9663 13887 9735
rect 14004 9663 14112 9735
rect 13776 6938 14112 9663
rect 13776 6866 13886 6938
rect 14003 6866 14112 6938
rect 13776 4392 14112 6866
rect 13776 4286 13830 4392
rect 13994 4286 14112 4392
rect 13776 4135 14112 4286
rect 13776 4060 13887 4135
rect 14000 4060 14112 4135
rect 13776 2440 14112 4060
rect 16464 22456 16800 22576
rect 16464 22400 16605 22456
rect 16661 22400 16800 22456
rect 16464 21769 16800 22400
rect 16464 21710 16593 21769
rect 16683 21710 16800 21769
rect 16464 20081 16800 21710
rect 16464 20022 16583 20081
rect 16673 20022 16800 20081
rect 16464 18969 16800 20022
rect 16464 18910 16593 18969
rect 16665 18910 16800 18969
rect 16464 18368 16800 18910
rect 16464 18258 16548 18368
rect 16719 18258 16800 18368
rect 16464 17278 16800 18258
rect 16464 17219 16599 17278
rect 16671 17219 16800 17278
rect 16464 16175 16800 17219
rect 16464 16114 16588 16175
rect 16667 16114 16800 16175
rect 16464 14478 16800 16114
rect 16464 14417 16592 14478
rect 16671 14417 16800 14478
rect 16464 13372 16800 14417
rect 16464 13308 16594 13372
rect 16668 13308 16800 13372
rect 16464 12809 16800 13308
rect 16464 12689 16544 12809
rect 16715 12689 16800 12809
rect 16464 11681 16800 12689
rect 16464 11617 16601 11681
rect 16675 11617 16800 11681
rect 16464 10574 16800 11617
rect 16464 10512 16593 10574
rect 16669 10512 16800 10574
rect 16464 8878 16800 10512
rect 16464 8816 16598 8878
rect 16674 8816 16800 8878
rect 16464 7772 16800 8816
rect 16464 7706 16589 7772
rect 16670 7706 16800 7772
rect 16464 7185 16800 7706
rect 16464 7065 16530 7185
rect 16701 7065 16800 7185
rect 16464 6082 16800 7065
rect 16464 6016 16593 6082
rect 16674 6016 16800 6082
rect 16464 4976 16800 6016
rect 16464 4906 16589 4976
rect 16672 4906 16800 4976
rect 16464 3288 16800 4906
rect 16464 3218 16594 3288
rect 16677 3218 16800 3288
rect 11648 2106 11758 2181
rect 11876 2106 11984 2181
rect 11648 1591 11984 2106
rect 11648 1471 11691 1591
rect 11862 1471 11984 1591
rect 11648 487 11984 1471
rect 11648 410 11760 487
rect 11872 410 11984 487
rect 11648 174 11984 410
rect 6778 -101 7112 0
rect 6778 -252 7113 -101
rect 6779 -745 7113 -252
rect 8570 -1002 8904 56
rect 11643 0 11984 174
rect 13775 1328 14114 2440
rect 13775 1255 13872 1328
rect 14002 1255 14114 1328
rect 11643 -252 11982 0
rect 11643 -748 11981 -252
rect 13775 -1002 14114 1255
rect 16464 2177 16800 3218
rect 16464 2104 16595 2177
rect 16675 2104 16800 2177
rect 16464 1596 16800 2104
rect 16464 1476 16552 1596
rect 16723 1476 16800 1596
rect 16464 485 16800 1476
rect 16464 412 16588 485
rect 16668 412 16800 485
rect 16464 56 16800 412
rect 16466 -252 16800 56
rect 18144 21179 18481 23184
rect 21284 22791 21631 28222
rect 23346 27247 23702 30202
rect 26155 28269 26502 28870
rect 26155 27940 26205 28269
rect 26457 27940 26502 28269
rect 18144 21103 18269 21179
rect 18354 21103 18481 21179
rect 18144 20943 18481 21103
rect 18144 20864 18268 20943
rect 18348 20864 18481 20943
rect 18144 18144 18481 20864
rect 18144 18065 18269 18144
rect 18349 18065 18481 18144
rect 18144 15598 18481 18065
rect 18144 15534 18260 15598
rect 18324 15534 18481 15598
rect 18144 15336 18481 15534
rect 18144 15261 18267 15336
rect 18351 15261 18481 15336
rect 18144 12530 18481 15261
rect 18144 12455 18268 12530
rect 18352 12455 18481 12530
rect 18144 9995 18481 12455
rect 18144 9896 18215 9995
rect 18370 9896 18481 9995
rect 18144 9735 18481 9896
rect 18144 9655 18265 9735
rect 18353 9655 18481 9735
rect 18144 6956 18481 9655
rect 18144 6876 18263 6956
rect 18351 6876 18481 6956
rect 18144 4397 18481 6876
rect 18144 4291 18225 4397
rect 18389 4291 18481 4397
rect 18144 4141 18481 4291
rect 18144 4066 18267 4141
rect 18360 4066 18481 4141
rect 18144 1335 18481 4066
rect 18144 1260 18262 1335
rect 18355 1260 18481 1335
rect 18144 123 18481 1260
rect 21280 22602 21631 22791
rect 23352 23240 23688 27247
rect 23352 23184 23493 23240
rect 23549 23184 23688 23240
rect 21280 22456 21616 22602
rect 21280 22400 21421 22456
rect 21477 22400 21616 22456
rect 21280 21773 21616 22400
rect 21280 21709 21412 21773
rect 21490 21709 21616 21773
rect 21280 20085 21616 21709
rect 21280 20021 21409 20085
rect 21486 20021 21616 20085
rect 21280 18978 21616 20021
rect 21280 18914 21404 18978
rect 21481 18914 21616 18978
rect 21280 18382 21616 18914
rect 21280 18262 21374 18382
rect 21545 18262 21616 18382
rect 21280 17285 21616 18262
rect 21280 17212 21407 17285
rect 21487 17212 21616 17285
rect 21280 16181 21616 17212
rect 21280 16108 21411 16181
rect 21491 16108 21616 16181
rect 21280 14481 21616 16108
rect 21280 14410 21397 14481
rect 21484 14410 21616 14481
rect 21280 13376 21616 14410
rect 21280 13305 21406 13376
rect 21493 13305 21616 13376
rect 21280 12819 21616 13305
rect 21280 12699 21367 12819
rect 21538 12699 21616 12819
rect 21280 11686 21616 12699
rect 21280 11610 21397 11686
rect 21483 11610 21616 11686
rect 21280 10576 21616 11610
rect 21280 10500 21402 10576
rect 21488 10500 21616 10576
rect 21280 8885 21616 10500
rect 21280 8811 21397 8885
rect 21484 8811 21616 8885
rect 21280 7779 21616 8811
rect 21280 7705 21404 7779
rect 21491 7705 21616 7779
rect 21280 7180 21616 7705
rect 21280 7060 21334 7180
rect 21505 7060 21616 7180
rect 21280 6083 21616 7060
rect 21280 6011 21400 6083
rect 21485 6011 21616 6083
rect 21280 4974 21616 6011
rect 21280 4902 21408 4974
rect 21493 4902 21616 4974
rect 21280 3283 21616 4902
rect 21280 3212 21401 3283
rect 21486 3212 21616 3283
rect 21280 2174 21616 3212
rect 21280 2103 21403 2174
rect 21488 2103 21616 2174
rect 21280 1576 21616 2103
rect 21280 1486 21377 1576
rect 21510 1486 21616 1576
rect 21280 480 21616 1486
rect 21280 408 21402 480
rect 21481 408 21616 480
rect 21280 198 21616 408
rect 16466 -717 16798 -252
rect 18144 -1002 18483 123
rect 21279 56 21616 198
rect 23352 21173 23688 23184
rect 26155 22632 26502 27940
rect 27780 27719 28136 30202
rect 23352 21097 23473 21173
rect 23558 21097 23688 21173
rect 23352 20944 23688 21097
rect 23352 20862 23462 20944
rect 23576 20862 23688 20944
rect 23352 18143 23688 20862
rect 23352 18068 23464 18143
rect 23575 18068 23688 18143
rect 23352 15598 23688 18068
rect 23352 15534 23473 15598
rect 23537 15534 23688 15598
rect 23352 15324 23688 15534
rect 23352 15258 23462 15324
rect 23577 15258 23688 15324
rect 23352 12526 23688 15258
rect 23352 12460 23462 12526
rect 23577 12460 23688 12526
rect 23352 9993 23688 12460
rect 23352 9894 23449 9993
rect 23604 9894 23688 9993
rect 23352 9726 23688 9894
rect 23352 9663 23463 9726
rect 23578 9663 23688 9726
rect 23352 6928 23688 9663
rect 23352 6865 23462 6928
rect 23577 6865 23688 6928
rect 23352 4397 23688 6865
rect 23352 4291 23429 4397
rect 23593 4291 23688 4397
rect 23352 4127 23688 4291
rect 23352 4056 23460 4127
rect 23576 4056 23688 4127
rect 23352 2343 23688 4056
rect 26152 22554 26502 22632
rect 27776 27380 28136 27719
rect 30972 28484 31319 29044
rect 30972 28204 31016 28484
rect 31278 28204 31319 28484
rect 27776 23251 28112 27380
rect 27776 23179 27862 23251
rect 28000 23179 28112 23251
rect 26152 22456 26488 22554
rect 26152 22400 26292 22456
rect 26348 22400 26488 22456
rect 26152 21776 26488 22400
rect 26152 21706 26264 21776
rect 26375 21706 26488 21776
rect 26152 20089 26488 21706
rect 26152 20017 26277 20089
rect 26366 20017 26488 20089
rect 26152 18975 26488 20017
rect 26152 18903 26281 18975
rect 26370 18903 26488 18975
rect 26152 18374 26488 18903
rect 26152 18254 26231 18374
rect 26402 18254 26488 18374
rect 26152 17285 26488 18254
rect 26152 17214 26270 17285
rect 26369 17214 26488 17285
rect 26152 16176 26488 17214
rect 26152 16105 26271 16176
rect 26370 16105 26488 16176
rect 26152 14483 26488 16105
rect 26152 14414 26265 14483
rect 26371 14414 26488 14483
rect 26152 13380 26488 14414
rect 26152 13311 26267 13380
rect 26373 13311 26488 13380
rect 26152 12819 26488 13311
rect 26152 12699 26218 12819
rect 26389 12699 26488 12819
rect 26152 11687 26488 12699
rect 26152 11611 26278 11687
rect 26367 11611 26488 11687
rect 26152 10582 26488 11611
rect 26152 10506 26277 10582
rect 26366 10506 26488 10582
rect 26152 8886 26488 10506
rect 26152 8811 26265 8886
rect 26364 8811 26488 8886
rect 26152 7783 26488 8811
rect 26152 7708 26273 7783
rect 26372 7708 26488 7783
rect 26152 7208 26488 7708
rect 26152 7088 26227 7208
rect 26398 7088 26488 7208
rect 26152 6090 26488 7088
rect 26152 6010 26275 6090
rect 26367 6010 26488 6090
rect 26152 4980 26488 6010
rect 26152 4900 26281 4980
rect 26373 4900 26488 4980
rect 26152 3290 26488 4900
rect 26152 3210 26264 3290
rect 26360 3210 26488 3290
rect 23352 1342 23690 2343
rect 23352 1271 23462 1342
rect 23578 1271 23690 1342
rect 21279 -252 21613 56
rect 23352 -252 23690 1271
rect 21281 -753 21610 -252
rect 23355 -1002 23690 -252
rect 26152 2179 26488 3210
rect 26152 2099 26276 2179
rect 26372 2099 26488 2179
rect 26152 1591 26488 2099
rect 26152 1471 26229 1591
rect 26400 1471 26488 1591
rect 26152 483 26488 1471
rect 26152 406 26275 483
rect 26363 406 26488 483
rect 26152 180 26488 406
rect 27776 21185 28112 23179
rect 30972 22874 31319 28204
rect 32923 26756 33279 30202
rect 35673 28867 36011 30202
rect 35672 28809 36011 28867
rect 40263 29131 40599 29343
rect 40263 29049 40384 29131
rect 40502 29049 40599 29131
rect 35672 27869 36008 28809
rect 40263 28012 40599 29049
rect 35672 27796 35784 27869
rect 35874 27796 36008 27869
rect 35672 26918 36008 27796
rect 35672 26846 35801 26918
rect 35890 26846 36008 26918
rect 27776 21109 27903 21185
rect 27988 21109 28112 21185
rect 27776 20937 28112 21109
rect 27776 20864 27887 20937
rect 28000 20864 28112 20937
rect 27776 18139 28112 20864
rect 27776 18066 27889 18139
rect 28002 18066 28112 18139
rect 27776 15600 28112 18066
rect 27776 15536 27903 15600
rect 27967 15536 28112 15600
rect 27776 12527 28112 15536
rect 27776 12456 27889 12527
rect 28001 12456 28112 12527
rect 27776 9981 28112 12456
rect 27776 9882 27863 9981
rect 28018 9882 28112 9981
rect 27776 9733 28112 9882
rect 27776 9663 27888 9733
rect 28000 9663 28112 9733
rect 27776 4397 28112 9663
rect 27776 4291 27849 4397
rect 28013 4291 28112 4397
rect 27776 4123 28112 4291
rect 27776 4050 27887 4123
rect 28001 4050 28112 4123
rect 27776 1330 28112 4050
rect 27776 1257 27887 1330
rect 28001 1257 28112 1330
rect 26152 -704 26491 180
rect 27776 -9 28112 1257
rect 30968 22728 31319 22874
rect 30968 22456 31304 22728
rect 30968 22400 31111 22456
rect 31167 22400 31304 22456
rect 30968 21771 31304 22400
rect 30968 21714 31080 21771
rect 31193 21714 31304 21771
rect 30968 20077 31304 21714
rect 30968 20020 31079 20077
rect 31192 20020 31304 20077
rect 30968 18969 31304 20020
rect 30968 18911 31080 18969
rect 31192 18911 31304 18969
rect 30968 18378 31304 18911
rect 30968 18258 31048 18378
rect 31219 18258 31304 18378
rect 30968 17279 31304 18258
rect 30968 17221 31080 17279
rect 31192 17221 31304 17279
rect 30968 16171 31304 17221
rect 30968 16115 31080 16171
rect 31192 16115 31304 16171
rect 30968 14479 31304 16115
rect 30968 14423 31080 14479
rect 31192 14423 31304 14479
rect 30968 13370 31304 14423
rect 30968 13310 31080 13370
rect 31192 13310 31304 13370
rect 30968 12814 31304 13310
rect 30968 12694 31032 12814
rect 31203 12694 31304 12814
rect 30968 11685 31304 12694
rect 30968 11625 31080 11685
rect 31192 11625 31304 11685
rect 30968 10574 31304 11625
rect 30968 10518 31080 10574
rect 31193 10518 31304 10574
rect 30968 8882 31304 10518
rect 30968 8826 31079 8882
rect 31192 8826 31304 8882
rect 30968 7772 31304 8826
rect 30968 7716 31079 7772
rect 31192 7716 31304 7772
rect 30968 7190 31304 7716
rect 30968 7070 31032 7190
rect 31203 7070 31304 7190
rect 30968 6082 31304 7070
rect 30968 6026 31080 6082
rect 31193 6026 31304 6082
rect 30968 4977 31304 6026
rect 30968 4921 31080 4977
rect 31192 4921 31304 4977
rect 30968 3278 31304 4921
rect 30968 3222 31080 3278
rect 31192 3222 31304 3278
rect 30968 2178 31304 3222
rect 30968 2117 31079 2178
rect 31193 2117 31304 2178
rect 30968 1595 31304 2117
rect 30968 1475 31033 1595
rect 31204 1475 31304 1595
rect 30968 482 31304 1475
rect 32928 21173 33264 26756
rect 32928 21097 33024 21173
rect 33109 21097 33264 21173
rect 32928 20938 33264 21097
rect 32928 20874 33039 20938
rect 33155 20874 33264 20938
rect 32928 18117 33264 20874
rect 32928 18053 33038 18117
rect 33154 18053 33264 18117
rect 32928 15605 33264 18053
rect 32928 15541 33057 15605
rect 33121 15541 33264 15605
rect 32928 15339 33264 15541
rect 32928 15269 33040 15339
rect 33152 15269 33264 15339
rect 32928 12535 33264 15269
rect 32928 12465 33040 12535
rect 33152 12465 33264 12535
rect 32928 9992 33264 12465
rect 32928 9893 33030 9992
rect 33185 9893 33264 9992
rect 32928 9732 33264 9893
rect 32928 9666 33031 9732
rect 33143 9666 33264 9732
rect 32928 6930 33264 9666
rect 32928 6864 33041 6930
rect 33153 6864 33264 6930
rect 32928 4392 33264 6864
rect 32928 4286 33020 4392
rect 33184 4286 33264 4392
rect 32928 4136 33264 4286
rect 32928 4072 33030 4136
rect 33139 4072 33264 4136
rect 32928 1329 33264 4072
rect 32928 1265 33043 1329
rect 33152 1265 33264 1329
rect 35672 25953 36008 26846
rect 37013 27079 37347 27150
rect 37013 27023 37124 27079
rect 37213 27023 37347 27079
rect 37013 26600 37347 27023
rect 37013 26314 37352 26600
rect 35672 25881 35794 25953
rect 35883 25881 36008 25953
rect 35672 24993 36008 25881
rect 35672 24915 35800 24993
rect 35893 24915 36008 24993
rect 35672 21175 36008 24915
rect 35672 21099 35797 21175
rect 35882 21099 36008 21175
rect 35672 20928 36008 21099
rect 35672 20869 35784 20928
rect 35896 20869 36008 20928
rect 35672 18127 36008 20869
rect 35672 18068 35784 18127
rect 35896 18068 36008 18127
rect 35672 15608 36008 18068
rect 35672 15544 35802 15608
rect 35866 15544 36008 15608
rect 35672 15333 36008 15544
rect 35672 15274 35784 15333
rect 35896 15274 36008 15333
rect 35672 12524 36008 15274
rect 35672 12465 35784 12524
rect 35896 12465 36008 12524
rect 35672 9981 36008 12465
rect 35672 9882 35753 9981
rect 35908 9882 36008 9981
rect 35672 9732 36008 9882
rect 35672 9674 35784 9732
rect 35896 9674 36008 9732
rect 35672 6921 36008 9674
rect 35672 6863 35784 6921
rect 35896 6863 36008 6921
rect 35672 4403 36008 6863
rect 35672 4297 35760 4403
rect 35924 4297 36008 4403
rect 35672 4130 36008 4297
rect 35672 4074 35783 4130
rect 35896 4074 36008 4130
rect 35672 1322 36008 4074
rect 32928 740 33264 1265
rect 30968 421 31079 482
rect 31193 421 31304 482
rect 30968 74 31304 421
rect 27776 -224 28113 -9
rect 27778 -1002 28113 -224
rect 30967 -112 31304 74
rect 32921 -56 33264 740
rect 35671 -56 36008 1322
rect 37016 26128 37352 26314
rect 37016 26063 37123 26128
rect 37244 26063 37352 26128
rect 37016 25163 37352 26063
rect 37016 25104 37126 25163
rect 37244 25104 37352 25163
rect 37016 24189 37352 25104
rect 37016 24130 37119 24189
rect 37237 24130 37352 24189
rect 37016 21773 37352 24130
rect 40262 22683 40600 24279
rect 37016 21707 37146 21773
rect 37224 21707 37352 21773
rect 37016 20089 37352 21707
rect 37016 20023 37145 20089
rect 37223 20023 37352 20089
rect 37016 18978 37352 20023
rect 37016 18909 37151 18978
rect 37227 18909 37352 18978
rect 37016 18374 37352 18909
rect 37016 18254 37093 18374
rect 37264 18254 37352 18374
rect 37016 17289 37352 18254
rect 37016 17220 37143 17289
rect 37219 17220 37352 17289
rect 37016 16175 37352 17220
rect 37016 16111 37144 16175
rect 37218 16111 37352 16175
rect 37016 14489 37352 16111
rect 37016 14425 37150 14489
rect 37224 14425 37352 14489
rect 37016 13376 37352 14425
rect 37016 13308 37148 13376
rect 37226 13308 37352 13376
rect 37016 12825 37352 13308
rect 37016 12705 37114 12825
rect 37285 12705 37352 12825
rect 37016 11686 37352 12705
rect 37016 11618 37146 11686
rect 37224 11618 37352 11686
rect 37016 10579 37352 11618
rect 37016 10506 37137 10579
rect 37219 10506 37352 10579
rect 37016 8885 37352 10506
rect 37016 8812 37142 8885
rect 37224 8812 37352 8885
rect 37016 7779 37352 8812
rect 37016 7711 37144 7779
rect 37228 7711 37352 7779
rect 37016 7194 37352 7711
rect 37016 7074 37088 7194
rect 37259 7074 37352 7194
rect 37016 6083 37352 7074
rect 37016 6015 37140 6083
rect 37224 6015 37352 6083
rect 37016 4976 37352 6015
rect 37016 4910 37140 4976
rect 37228 4910 37352 4976
rect 37016 3285 37352 4910
rect 37016 3219 37137 3285
rect 37225 3219 37352 3285
rect 37016 1597 37352 3219
rect 37016 1477 37103 1597
rect 37274 1477 37352 1597
rect 37016 -56 37352 1477
rect 30967 -252 31301 -112
rect 30967 -754 31300 -252
rect -2581 -1006 28113 -1002
rect 32921 -1006 33262 -56
rect 35671 -1006 36007 -56
rect 37018 -252 37352 -56
rect 37019 -775 37350 -252
rect 44357 -1006 47058 30202
rect -2581 -1009 47058 -1006
rect -6233 -1012 47058 -1009
rect -6233 -3603 47061 -1012
rect 44357 -3640 47058 -3603
use 4MSB_weighted_binary  4MSB_weighted_binary_0
timestamp 1755923935
transform -1 0 43959 0 1 27999
box 2352 -4032 10080 56
use 6MSB_MATRIX  6MSB_MATRIX_0
timestamp 1755923713
transform 1 0 -2298 0 1 21392
box 2298 -21392 43904 2632
<< labels >>
flabel metal2 25302 39863 26122 40690 1 FreeSans 8000 0 0 0 X5
port 5 n
flabel metal2 21605 39810 22425 40637 1 FreeSans 8000 0 0 0 X7
port 7 n
flabel metal2 11162 39568 11982 39838 1 FreeSans 8000 0 0 0 X8
port 8 n
flabel metal2 8115 39645 8935 40472 1 FreeSans 8000 0 0 0 X10
port 10 n
flabel metal2 34952 39984 35772 40811 1 FreeSans 8000 0 0 0 X1
port 1 n
flabel metal2 32703 39616 33523 40447 1 FreeSans 8000 0 0 0 X2
port 2 n
flabel metal2 36320 39983 37140 40814 1 FreeSans 6400 0 0 0 X4
port 4 n
flabel metal2 31082 40348 31902 41179 1 FreeSans 6400 0 0 0 X3
port 3 n
flabel space 38229 38817 39049 39648 1 FreeSans 8000 0 0 0 CLK
port 11 n
flabel metal2 3166 39659 3986 40486 1 FreeSans 8000 0 0 0 X9
port 9 n
flabel metal2 16947 39645 17767 40472 1 FreeSans 8000 0 0 0 X6
port 6 n
flabel metal2 52171 30107 53635 31531 1 FreeSans 8000 0 0 0 VBIAS
port 14 n
flabel metal2 55903 27782 57367 29206 1 FreeSans 8000 0 0 0 OUTP
port 12 n
flabel space 53438 24944 54902 26369 1 FreeSans 8000 0 0 0 OUTN
port 13 n
flabel metal4 -6208 30202 46994 32676 1 FreeSans 11200 0 0 0 VDD
port 15 n
flabel metal3 -10148 34395 50919 36995 1 FreeSans 11200 0 0 0 VSS
port 16 n
flabel metal3 48434 -7526 50908 37079 1 FreeSans 11200 0 0 0 VSS
port 16 n
flabel metal3 -10147 -7526 50920 -4926 1 FreeSans 11200 0 0 0 VSS
port 16 n
flabel metal3 -10148 -7521 -7674 37008 1 FreeSans 11200 0 0 0 VSS
port 16 n
flabel metal4 -6233 -3603 47061 -1012 1 FreeSans 11200 0 0 0 VDD
port 15 n
flabel metal4 44357 -3640 47058 30206 1 FreeSans 11200 0 0 0 VDD
port 15 n
flabel metal4 -6233 -3603 -3581 30269 1 FreeSans 11200 0 0 0 VDD
port 15 n
<< end >>
