magic
tech gf180mcuD
magscale 1 10
timestamp 1754367086
<< pwell >>
rect 519 1024 1664 1719
<< nmos >>
rect 728 1400 784 1444
rect 956 1400 1012 1444
rect 1292 1366 1348 1478
rect 1440 1360 1500 1484
<< ndiff >>
rect 602 1446 682 1462
rect 602 1398 618 1446
rect 666 1444 682 1446
rect 830 1446 910 1462
rect 830 1444 846 1446
rect 666 1400 728 1444
rect 784 1400 846 1444
rect 666 1398 682 1400
rect 602 1382 682 1398
rect 830 1398 846 1400
rect 894 1444 910 1446
rect 1394 1478 1440 1484
rect 1246 1462 1292 1478
rect 1058 1446 1138 1462
rect 1058 1444 1074 1446
rect 894 1400 956 1444
rect 1012 1400 1074 1444
rect 894 1398 910 1400
rect 830 1382 910 1398
rect 1058 1398 1074 1400
rect 1122 1398 1138 1446
rect 1058 1382 1138 1398
rect 1198 1446 1292 1462
rect 1198 1398 1214 1446
rect 1262 1398 1292 1446
rect 1198 1382 1292 1398
rect 1246 1366 1292 1382
rect 1348 1366 1440 1478
rect 1394 1360 1440 1366
rect 1500 1462 1546 1484
rect 1500 1446 1596 1462
rect 1500 1398 1532 1446
rect 1580 1398 1596 1446
rect 1500 1382 1596 1398
rect 1500 1360 1546 1382
<< ndiffc >>
rect 618 1398 666 1446
rect 846 1398 894 1446
rect 1074 1398 1122 1446
rect 1214 1398 1262 1446
rect 1532 1398 1580 1446
<< polysilicon >>
rect 716 1554 796 1570
rect 716 1506 732 1554
rect 780 1506 796 1554
rect 716 1490 796 1506
rect 944 1554 1024 1570
rect 944 1506 960 1554
rect 1008 1506 1024 1554
rect 944 1490 1024 1506
rect 1292 1568 1500 1581
rect 1292 1522 1350 1568
rect 1450 1522 1500 1568
rect 1292 1504 1500 1522
rect 728 1444 784 1490
rect 728 1354 784 1400
rect 956 1444 1012 1490
rect 1292 1478 1348 1504
rect 1440 1484 1500 1504
rect 956 1354 1012 1400
rect 1292 1320 1348 1366
rect 1440 1314 1500 1360
<< polycontact >>
rect 732 1506 780 1554
rect 960 1506 1008 1554
rect 1350 1522 1450 1568
<< metal1 >>
rect 612 1460 672 1588
rect 726 1554 786 1628
rect 726 1506 732 1554
rect 780 1506 786 1554
rect 726 1494 786 1506
rect 954 1554 1014 1632
rect 954 1506 960 1554
rect 1008 1506 1014 1554
rect 954 1494 1014 1506
rect 1068 1460 1128 1588
rect 1315 1568 1478 1576
rect 1315 1522 1350 1568
rect 1450 1522 1478 1568
rect 1315 1512 1478 1522
rect 604 1446 680 1460
rect 604 1398 618 1446
rect 666 1398 680 1446
rect 604 1384 680 1398
rect 832 1446 908 1460
rect 832 1398 846 1446
rect 894 1398 908 1446
rect 832 1384 908 1398
rect 1060 1446 1136 1460
rect 1060 1398 1074 1446
rect 1122 1398 1136 1446
rect 1060 1384 1136 1398
rect 1200 1446 1276 1460
rect 1200 1398 1214 1446
rect 1262 1398 1276 1446
rect 1200 1384 1276 1398
rect 1518 1446 1594 1460
rect 1518 1398 1532 1446
rect 1580 1398 1594 1446
rect 1518 1384 1594 1398
rect 846 1332 894 1384
rect 1214 1332 1262 1384
rect 846 1284 1262 1332
rect 1152 1283 1262 1284
rect 1532 1231 1580 1384
rect 604 1120 1624 1231
<< labels >>
flabel metal1 726 1494 786 1628 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 954 1494 1014 1632 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 612 1392 672 1588 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 1068 1392 1128 1588 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 1315 1512 1478 1576 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel pwell 619 1123 734 1226 1 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
flabel metal1 784 1120 1624 1231 1 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional
<< end >>
