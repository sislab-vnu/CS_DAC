magic
tech gf180mcuD
magscale 1 10
timestamp 1756789507
<< isosubstrate >>
rect 6892 942 6906 1152
rect 7492 966 7548 1130
rect 6892 860 6904 942
rect 6892 504 6904 757
<< pwell >>
rect 6892 942 6906 1152
rect 7492 966 7548 1130
rect 6892 860 6904 942
rect 6892 504 6904 757
rect 7112 -216 7168 44
rect 7214 -125 7242 -81
rect 6805 -590 7966 -456
rect 8232 -1176 8288 -1120
rect 6804 -1710 8212 -1575
rect 6892 -2344 6964 -2161
rect 6892 -2407 7096 -2344
rect 7485 -2378 7541 -2184
rect 6893 -2595 7096 -2407
rect 6890 -2603 7096 -2595
rect 6890 -2649 6968 -2603
rect 6805 -2830 8325 -2649
rect 6890 -2856 6968 -2830
<< psubdiff >>
rect 2672 623 2772 640
rect 2672 557 2691 623
rect 2751 557 2772 623
rect 2672 540 2772 557
rect 2672 -503 2772 -480
rect 2672 -560 2692 -503
rect 2748 -560 2772 -503
rect 2672 -580 2772 -560
rect 2672 -1622 2772 -1600
rect 2672 -1682 2694 -1622
rect 2753 -1682 2772 -1622
rect 2672 -1700 2772 -1682
rect 2672 -2736 2772 -2720
rect 2672 -2800 2689 -2736
rect 2750 -2800 2772 -2736
rect 2672 -2820 2772 -2800
<< nsubdiff >>
rect 2672 1407 2772 1424
rect 2672 1341 2690 1407
rect 2750 1341 2772 1407
rect 2672 1324 2772 1341
rect 2672 280 2772 304
rect 2672 223 2693 280
rect 2749 223 2772 280
rect 2672 204 2772 223
rect 2672 -840 2772 -816
rect 2672 -900 2691 -840
rect 2750 -900 2772 -840
rect 2672 -916 2772 -900
rect 2672 -1956 2772 -1936
rect 2672 -2020 2691 -1956
rect 2752 -2020 2772 -1956
rect 2672 -2036 2772 -2020
<< psubdiffcont >>
rect 2691 557 2751 623
rect 2692 -560 2748 -503
rect 2694 -1682 2753 -1622
rect 2689 -2800 2750 -2736
<< nsubdiffcont >>
rect 2690 1341 2750 1407
rect 2693 223 2749 280
rect 2691 -900 2750 -840
rect 2691 -2020 2752 -1956
<< metal1 >>
rect 2128 1020 2464 1680
rect 7085 1400 8214 1456
rect 8270 1400 8288 1456
rect 2128 944 2801 1020
rect 5936 952 6273 1008
rect 2128 -100 2464 944
rect 7085 882 7141 1400
rect 8456 1288 8792 1624
rect 7492 1232 8792 1288
rect 7492 882 7548 1232
rect 7668 1064 8220 1120
rect 8276 1064 8288 1120
rect 6806 530 7923 682
rect 7112 280 8211 336
rect 8267 280 8288 336
rect 2128 -176 2803 -100
rect 5936 -139 6324 -112
rect 5944 -168 6260 -139
rect 2128 -1220 2464 -176
rect 7112 -216 7168 280
rect 8456 168 8792 1232
rect 7516 112 8792 168
rect 7516 -216 7572 112
rect 7694 -56 8220 0
rect 8276 -56 8288 0
rect 6805 -590 7966 -456
rect 7367 -840 8216 -784
rect 8272 -840 8288 -784
rect 2128 -1296 2802 -1220
rect 5929 -1288 6277 -1232
rect 2128 -2340 2464 -1296
rect 7367 -1327 7423 -840
rect 8456 -952 8792 112
rect 7784 -1008 8792 -952
rect 7784 -1327 7840 -1008
rect 7956 -1176 8218 -1120
rect 8274 -1176 8288 -1120
rect 6804 -1710 8212 -1575
rect 7112 -1960 8217 -1904
rect 8273 -1960 8288 -1904
rect 2128 -2352 2804 -2340
rect 2128 -2408 2806 -2352
rect 5936 -2407 6272 -2352
rect 2128 -2416 2804 -2408
rect 2128 -2968 2464 -2416
rect 7112 -2496 7168 -1960
rect 8456 -2072 8792 -1008
rect 7616 -2128 8792 -2072
rect 7616 -2496 7672 -2128
rect 7844 -2352 8275 -2296
rect 8331 -2352 8344 -2296
rect 6805 -2830 8325 -2649
rect 8456 -2912 8792 -2128
rect 8960 1456 9296 1624
rect 8960 1400 9072 1456
rect 9184 1400 9296 1456
rect 8960 336 9296 1400
rect 8960 280 9072 336
rect 9184 280 9296 336
rect 8960 -784 9296 280
rect 8960 -840 9072 -784
rect 9184 -840 9296 -784
rect 8960 -1904 9296 -840
rect 8960 -1960 9072 -1904
rect 9184 -1960 9296 -1904
rect 8960 -2912 9296 -1960
rect 9464 1120 9800 1624
rect 9464 1064 9576 1120
rect 9688 1064 9800 1120
rect 9464 0 9800 1064
rect 9464 -56 9576 0
rect 9688 -56 9800 0
rect 9464 -1120 9800 -56
rect 9464 -1176 9576 -1120
rect 9688 -1176 9800 -1120
rect 9464 -2296 9800 -1176
rect 9464 -2352 9576 -2296
rect 9688 -2352 9800 -2296
rect 9464 -2912 9800 -2352
<< via1 >>
rect 8214 1400 8270 1456
rect 5432 1344 5544 1400
rect 6397 1176 6453 1232
rect 6496 952 6552 1008
rect 3583 850 3639 906
rect 7206 1017 7262 1073
rect 7374 1017 7430 1073
rect 8220 1064 8276 1120
rect 3808 560 3920 616
rect 8211 280 8267 336
rect 5432 224 5544 280
rect 6396 56 6452 112
rect 6496 -179 6552 -123
rect 3582 -271 3638 -215
rect 7224 -84 7280 -28
rect 7400 -83 7456 -27
rect 8220 -56 8276 0
rect 3808 -560 3920 -504
rect 8216 -840 8272 -784
rect 5432 -896 5544 -840
rect 6398 -1064 6454 -1008
rect 6496 -1288 6552 -1232
rect 7487 -1195 7543 -1139
rect 7662 -1195 7718 -1139
rect 8218 -1176 8274 -1120
rect 3583 -1390 3639 -1334
rect 3808 -1680 3920 -1624
rect 8217 -1960 8273 -1904
rect 5432 -2016 5544 -1960
rect 6395 -2240 6451 -2184
rect 6496 -2408 6552 -2352
rect 3583 -2511 3639 -2455
rect 7257 -2376 7313 -2320
rect 7485 -2378 7541 -2322
rect 8275 -2352 8331 -2296
rect 3808 -2800 3920 -2744
rect 9072 1400 9184 1456
rect 9072 280 9184 336
rect 9072 -840 9184 -784
rect 9072 -1960 9184 -1904
rect 9576 1064 9688 1120
rect 9576 -56 9688 0
rect 9576 -1176 9688 -1120
rect 9576 -2352 9688 -2296
<< metal2 >>
rect 8198 1456 8285 1467
rect 9044 1456 9211 1482
rect 5417 1400 5557 1412
rect 5417 1344 5432 1400
rect 5544 1344 5557 1400
rect 8198 1400 8214 1456
rect 8270 1400 9072 1456
rect 9184 1400 9240 1456
rect 8198 1384 8285 1400
rect 9044 1367 9211 1400
rect 5417 1332 5557 1344
rect 6387 1232 6463 1242
rect 6387 1176 6397 1232
rect 6453 1176 7430 1232
rect 6387 1166 6463 1176
rect 3576 906 3657 1132
rect 7374 1082 7430 1176
rect 8205 1120 8288 1137
rect 9551 1120 9716 1147
rect 7196 1073 7272 1082
rect 7196 1017 7206 1073
rect 7262 1017 7272 1073
rect 6478 1008 6564 1014
rect 7196 1008 7272 1017
rect 6478 952 6496 1008
rect 6552 952 7272 1008
rect 7364 1073 7440 1082
rect 7364 1017 7374 1073
rect 7430 1017 7440 1073
rect 8205 1064 8220 1120
rect 8276 1064 9576 1120
rect 9688 1064 9744 1120
rect 8205 1048 8288 1064
rect 9551 1041 9716 1064
rect 7364 1006 7440 1017
rect 6478 931 6564 952
rect 3576 850 3583 906
rect 3639 850 3657 906
rect 3576 832 3657 850
rect 3798 616 3934 627
rect 3798 560 3808 616
rect 3920 560 3934 616
rect 3798 550 3934 560
rect 8195 336 8278 355
rect 9042 336 9211 363
rect 5417 280 5558 291
rect 5417 224 5432 280
rect 5544 224 5558 280
rect 8195 280 8211 336
rect 8267 280 9072 336
rect 9184 280 9240 336
rect 8195 263 8278 280
rect 9042 250 9211 280
rect 5417 213 5558 224
rect 6384 112 6460 122
rect 6384 56 6396 112
rect 6452 56 7456 112
rect 6384 46 6460 56
rect 3576 -215 3657 12
rect 7400 -18 7456 56
rect 8203 0 8288 14
rect 9544 0 9713 27
rect 7214 -28 7290 -18
rect 7214 -84 7224 -28
rect 7280 -84 7290 -28
rect 7214 -94 7290 -84
rect 7390 -27 7466 -18
rect 7390 -83 7400 -27
rect 7456 -83 7466 -27
rect 8203 -56 8220 0
rect 8276 -56 9576 0
rect 9688 -56 9744 0
rect 8203 -69 8288 -56
rect 9544 -82 9713 -56
rect 7390 -94 7466 -83
rect 6481 -123 6564 -106
rect 7214 -123 7280 -94
rect 6481 -179 6496 -123
rect 6552 -179 7280 -123
rect 6481 -189 6564 -179
rect 3576 -271 3582 -215
rect 3638 -271 3657 -215
rect 3576 -288 3657 -271
rect 3796 -504 3932 -494
rect 3796 -560 3808 -504
rect 3920 -560 3932 -504
rect 3796 -575 3932 -560
rect 8196 -784 8288 -761
rect 9042 -784 9214 -754
rect 5421 -840 5555 -832
rect 5421 -896 5432 -840
rect 5544 -896 5555 -840
rect 8196 -840 8216 -784
rect 8272 -840 9072 -784
rect 9184 -840 9240 -784
rect 8196 -861 8288 -840
rect 9042 -869 9214 -840
rect 5421 -910 5555 -896
rect 6387 -1008 6468 -1000
rect 6387 -1064 6398 -1008
rect 6454 -1064 7718 -1008
rect 6387 -1073 6468 -1064
rect 3576 -1334 3657 -1108
rect 7662 -1129 7718 -1064
rect 8206 -1120 8282 -1109
rect 9547 -1120 9719 -1090
rect 7476 -1139 7552 -1129
rect 7476 -1195 7487 -1139
rect 7543 -1195 7552 -1139
rect 6482 -1232 6564 -1226
rect 7476 -1232 7552 -1195
rect 7652 -1139 7728 -1129
rect 7652 -1195 7662 -1139
rect 7718 -1195 7728 -1139
rect 8206 -1176 8218 -1120
rect 8274 -1176 9576 -1120
rect 9688 -1176 9744 -1120
rect 8206 -1185 8282 -1176
rect 7652 -1205 7728 -1195
rect 9547 -1207 9719 -1176
rect 6482 -1288 6496 -1232
rect 6552 -1288 7552 -1232
rect 6482 -1309 6564 -1288
rect 3576 -1390 3583 -1334
rect 3639 -1390 3657 -1334
rect 3576 -1408 3657 -1390
rect 3796 -1624 3932 -1613
rect 3796 -1680 3808 -1624
rect 3920 -1680 3932 -1624
rect 3796 -1691 3932 -1680
rect 8201 -1904 8288 -1889
rect 9045 -1904 9208 -1881
rect 5421 -1960 5554 -1950
rect 5421 -2016 5432 -1960
rect 5544 -2016 5554 -1960
rect 8201 -1960 8217 -1904
rect 8273 -1960 9072 -1904
rect 9184 -1960 9240 -1904
rect 8201 -1974 8288 -1960
rect 9045 -1987 9208 -1960
rect 5421 -2027 5554 -2016
rect 6384 -2184 6460 -2174
rect 3576 -2455 3657 -2228
rect 6384 -2240 6395 -2184
rect 6451 -2240 7541 -2184
rect 6384 -2250 6460 -2240
rect 7485 -2312 7541 -2240
rect 8264 -2296 8340 -2286
rect 9547 -2296 9716 -2268
rect 7247 -2320 7323 -2312
rect 6483 -2352 6564 -2346
rect 7247 -2352 7257 -2320
rect 6483 -2408 6496 -2352
rect 6552 -2376 7257 -2352
rect 7313 -2376 7323 -2320
rect 6552 -2408 7323 -2376
rect 7475 -2322 7551 -2312
rect 7475 -2378 7485 -2322
rect 7541 -2378 7551 -2322
rect 8264 -2352 8275 -2296
rect 8331 -2352 9576 -2296
rect 9688 -2352 9744 -2296
rect 8264 -2362 8340 -2352
rect 7475 -2388 7551 -2378
rect 9547 -2381 9716 -2352
rect 6483 -2429 6564 -2408
rect 3576 -2511 3583 -2455
rect 3639 -2511 3657 -2455
rect 3576 -2528 3657 -2511
rect 3795 -2744 3934 -2731
rect 3795 -2800 3808 -2744
rect 3920 -2800 3934 -2744
rect 3795 -2811 3934 -2800
<< via2 >>
rect 5432 1344 5544 1400
rect 3808 560 3920 616
rect 5432 224 5544 280
rect 3808 -560 3920 -504
rect 5432 -896 5544 -840
rect 3808 -1680 3920 -1624
rect 5432 -2016 5544 -1960
rect 3808 -2800 3920 -2744
<< metal3 >>
rect 3751 616 3977 1678
rect 3751 560 3808 616
rect 3920 560 3977 616
rect 3751 -504 3977 560
rect 3751 -560 3808 -504
rect 3920 -560 3977 -504
rect 3751 -1624 3977 -560
rect 3751 -1680 3808 -1624
rect 3920 -1680 3977 -1624
rect 3751 -2744 3977 -1680
rect 3751 -2800 3808 -2744
rect 3920 -2800 3977 -2744
rect 3751 -3026 3977 -2800
rect 5376 1400 5600 1680
rect 5376 1344 5432 1400
rect 5544 1344 5600 1400
rect 5376 280 5600 1344
rect 5376 224 5432 280
rect 5544 224 5600 280
rect 5376 -840 5600 224
rect 5376 -896 5432 -840
rect 5544 -896 5600 -840
rect 5376 -1960 5600 -896
rect 5376 -2016 5432 -1960
rect 5544 -2016 5600 -1960
rect 5376 -3024 5600 -2016
use CS_Switch_1x1  CS_Switch_1x1_0
timestamp 1755764817
transform 1 0 7206 0 1 938
box -306 -434 837 214
use CS_Switch_2x2  CS_Switch_2x2_1
timestamp 1755705199
transform 1 0 7248 0 1 -180
box -356 -436 795 224
use CS_Switch_4x2  CS_Switch_4x2_0
timestamp 1755705775
transform 1 0 7196 0 1 -1551
box -304 -185 1117 488
use CS_Switch_8x2  CS_Switch_8x2_0
timestamp 1755706082
transform 1 0 6529 0 1 -3880
box 426 1024 1804 1719
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2662 0 1 -2770
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_1
timestamp 1753044640
transform 1 0 2662 0 1 590
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_2
timestamp 1753044640
transform 1 0 2662 0 1 -530
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_3
timestamp 1753044640
transform 1 0 2662 0 1 -1650
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 6134 0 1 -530
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_1
timestamp 1753044640
transform 1 0 6134 0 1 590
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_2
timestamp 1753044640
transform 1 0 6134 0 1 -2770
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_3
timestamp 1753044640
transform 1 0 6134 0 1 -1650
box -86 -86 758 870
<< labels >>
flabel metal1 9464 -2912 9800 1624 1 FreeSans 800 0 0 0 VBIAS
port 7 n
flabel metal1 8456 -2912 8792 1624 1 FreeSans 800 0 0 0 OUTN
port 6 n
flabel metal1 8960 -2912 9296 1624 1 FreeSans 800 0 0 0 OUTP
port 5 n
flabel metal2 3576 832 3657 1132 1 FreeSans 800 0 0 0 D1
port 1 n
flabel metal2 3576 -288 3657 12 1 FreeSans 800 0 0 0 D2
port 2 n
flabel metal2 3576 -1408 3657 -1108 1 FreeSans 800 0 0 0 D3
port 3 n
flabel metal2 3576 -2528 3657 -2228 1 FreeSans 800 0 0 0 D4
port 4 n
flabel metal1 2128 -2968 2464 1680 1 FreeSans 800 0 0 0 CLK
port 8 n
flabel metal3 5376 -3024 5600 1680 1 FreeSans 800 0 0 0 VDD
port 9 n
flabel metal3 3751 -3026 3977 1678 1 FreeSans 800 0 0 0 VSS
port 10 n
<< properties >>
string CS_Switch_2x2_0 x1
string name x1
<< end >>
