magic
tech gf180mcuD
magscale 1 10
timestamp 1758595292
<< metal1 >>
rect 40152 41384 40488 42000
rect 40824 41664 91560 41720
rect 40824 41640 42392 41664
rect 40824 41584 41188 41640
rect 41244 41584 42392 41640
rect 40824 41552 42392 41584
rect 42504 41552 43756 41664
rect 43868 41552 45212 41664
rect 45324 41640 48720 41664
rect 45324 41584 47516 41640
rect 47572 41584 48720 41640
rect 45324 41552 48720 41584
rect 48832 41552 50088 41664
rect 50200 41552 51550 41664
rect 51662 41640 55048 41664
rect 51662 41584 53844 41640
rect 53900 41584 55048 41640
rect 51662 41552 55048 41584
rect 55160 41552 56416 41664
rect 56528 41552 57873 41664
rect 57985 41640 61376 41664
rect 57985 41584 60172 41640
rect 60228 41584 61376 41640
rect 57985 41552 61376 41584
rect 61488 41552 62746 41664
rect 62858 41552 64204 41664
rect 64316 41640 67704 41664
rect 64316 41584 66500 41640
rect 66556 41584 67704 41640
rect 64316 41552 67704 41584
rect 67816 41552 69077 41664
rect 69189 41552 70528 41664
rect 70640 41640 74032 41664
rect 70640 41584 72828 41640
rect 72884 41584 74032 41640
rect 70640 41552 74032 41584
rect 74144 41552 75403 41664
rect 75515 41552 76860 41664
rect 76972 41640 80360 41664
rect 76972 41584 79156 41640
rect 79212 41584 80360 41640
rect 76972 41552 80360 41584
rect 80472 41552 81734 41664
rect 81846 41552 83186 41664
rect 83298 41642 91560 41664
rect 83298 41584 85231 41642
rect 85288 41584 91560 41642
rect 83298 41552 91560 41584
rect 40824 41496 91560 41552
rect 40152 41300 91560 41384
rect 40152 41244 41357 41300
rect 41413 41244 47685 41300
rect 47741 41244 54013 41300
rect 54069 41244 60341 41300
rect 60397 41244 66669 41300
rect 66725 41244 72997 41300
rect 73053 41244 79325 41300
rect 79381 41244 91560 41300
rect 40152 41160 91560 41244
rect 40152 37800 40488 41160
rect 40824 40992 91560 41048
rect 40824 40965 91363 40992
rect 40824 40909 46844 40965
rect 46900 40909 53172 40965
rect 53228 40909 59500 40965
rect 59556 40909 65828 40965
rect 65884 40909 72156 40965
rect 72212 40909 78484 40965
rect 78540 40909 84812 40965
rect 84868 40909 91363 40965
rect 40824 40880 91363 40909
rect 91475 40880 91560 40992
rect 40824 40824 91560 40880
rect 91672 40712 92008 42056
rect 40824 40489 92008 40712
rect 40824 40488 85344 40489
rect 91350 40488 92008 40489
rect 41160 40405 41272 40432
rect 41160 40349 41189 40405
rect 41245 40349 41272 40405
rect 41160 39144 41272 40349
rect 41328 40405 41440 40432
rect 41328 40349 41363 40405
rect 41419 40349 41440 40405
rect 41328 39980 41440 40349
rect 41328 39904 41709 39980
rect 46348 39802 46424 40488
rect 46816 40405 46928 40432
rect 46816 40349 46844 40405
rect 46900 40349 46928 40405
rect 46816 40320 46928 40349
rect 47488 40400 47600 40432
rect 47488 40344 47517 40400
rect 47573 40344 47600 40400
rect 46830 39802 46906 40320
rect 47488 39144 47600 40344
rect 47656 40405 47768 40432
rect 47656 40349 47685 40405
rect 47741 40349 47768 40405
rect 47656 39980 47768 40349
rect 47656 39904 48037 39980
rect 52676 39802 52752 40488
rect 53144 40405 53256 40432
rect 53144 40349 53172 40405
rect 53228 40349 53256 40405
rect 53144 40320 53256 40349
rect 53816 40404 53928 40432
rect 53816 40348 53841 40404
rect 53897 40348 53928 40404
rect 53158 39802 53234 40320
rect 53816 39144 53928 40348
rect 53984 40405 54096 40432
rect 53984 40349 54016 40405
rect 54072 40349 54096 40405
rect 53984 39980 54096 40349
rect 53984 39904 54365 39980
rect 59004 39802 59080 40488
rect 59472 40405 59584 40432
rect 59472 40349 59500 40405
rect 59556 40349 59584 40405
rect 59472 40320 59584 40349
rect 60144 40406 60256 40432
rect 60144 40350 60173 40406
rect 60229 40350 60256 40406
rect 59486 39802 59562 40320
rect 60144 39144 60256 40350
rect 60312 40403 60424 40432
rect 60312 40347 60344 40403
rect 60400 40347 60424 40403
rect 60312 39980 60424 40347
rect 60312 39904 60693 39980
rect 65332 39802 65408 40488
rect 65800 40405 65912 40432
rect 65800 40349 65828 40405
rect 65884 40349 65912 40405
rect 65800 40320 65912 40349
rect 66472 40405 66584 40432
rect 66472 40349 66501 40405
rect 66557 40349 66584 40405
rect 65814 39802 65890 40320
rect 66472 39144 66584 40349
rect 66640 40405 66752 40432
rect 66640 40349 66673 40405
rect 66729 40349 66752 40405
rect 66640 39980 66752 40349
rect 66640 39904 67021 39980
rect 71660 39802 71736 40488
rect 72128 40405 72240 40432
rect 72128 40349 72156 40405
rect 72212 40349 72240 40405
rect 72128 40320 72240 40349
rect 72800 40405 72912 40432
rect 72800 40349 72829 40405
rect 72885 40349 72912 40405
rect 72142 39802 72218 40320
rect 72800 39144 72912 40349
rect 72968 40403 73080 40432
rect 72968 40347 72997 40403
rect 73053 40347 73080 40403
rect 72968 39980 73080 40347
rect 72968 39904 73349 39980
rect 77988 39802 78064 40488
rect 78456 40405 78568 40432
rect 78456 40349 78484 40405
rect 78540 40349 78568 40405
rect 78456 40320 78568 40349
rect 79128 40403 79240 40432
rect 79128 40347 79158 40403
rect 79214 40347 79240 40403
rect 78470 39802 78546 40320
rect 79128 39144 79240 40347
rect 79296 40400 79408 40432
rect 79296 40344 79328 40400
rect 79384 40344 79408 40400
rect 79296 39980 79408 40344
rect 79296 39904 79677 39980
rect 84316 39802 84392 40488
rect 84784 40405 84896 40432
rect 84784 40349 84812 40405
rect 84868 40349 84896 40405
rect 84784 40320 84896 40349
rect 84798 39802 84874 40320
rect 41160 39032 41749 39144
rect 47488 39032 48077 39144
rect 53816 39032 54405 39144
rect 60144 39032 60733 39144
rect 66472 39032 67061 39144
rect 72800 39032 73389 39144
rect 79128 39032 79717 39144
rect 40824 38416 91560 38472
rect 40824 38386 91363 38416
rect 40824 38330 46811 38386
rect 46867 38330 53139 38386
rect 53195 38330 59467 38386
rect 59523 38330 65795 38386
rect 65851 38330 72123 38386
rect 72179 38330 78451 38386
rect 78507 38330 84779 38386
rect 84835 38330 91363 38386
rect 40824 38304 91363 38330
rect 91475 38304 91560 38416
rect 40824 38248 91560 38304
rect 40544 38080 91560 38136
rect 40544 37968 40626 38080
rect 40738 38056 91560 38080
rect 40738 38000 41188 38056
rect 41244 38053 47516 38056
rect 41244 38000 43429 38053
rect 40738 37997 43429 38000
rect 43485 38000 47516 38053
rect 47572 38053 53844 38056
rect 47572 38000 49757 38053
rect 43485 37997 49757 38000
rect 49813 38000 53844 38053
rect 53900 38053 60172 38056
rect 53900 38000 56085 38053
rect 49813 37997 56085 38000
rect 56141 38000 60172 38053
rect 60228 38053 66500 38056
rect 60228 38000 62413 38053
rect 56141 37997 62413 38000
rect 62469 38000 66500 38053
rect 66556 38053 72828 38056
rect 66556 38000 68741 38053
rect 62469 37997 68741 38000
rect 68797 38000 72828 38053
rect 72884 38053 79156 38056
rect 72884 38000 75069 38053
rect 68797 37997 75069 38000
rect 75125 38000 79156 38053
rect 79212 38053 85484 38056
rect 79212 38000 81397 38053
rect 75125 37997 81397 38000
rect 81453 38000 85484 38053
rect 85540 38000 91560 38056
rect 81453 37997 91560 38000
rect 40738 37968 91560 37997
rect 40544 37912 91560 37968
rect 40152 37716 91560 37800
rect 40152 37660 41357 37716
rect 41413 37660 47685 37716
rect 47741 37660 54013 37716
rect 54069 37660 60341 37716
rect 60397 37660 66669 37716
rect 66725 37660 72997 37716
rect 73053 37660 79325 37716
rect 79381 37660 85653 37716
rect 85709 37660 91560 37716
rect 40152 37576 91560 37660
rect 40152 34216 40488 37576
rect 40824 37408 91560 37464
rect 40824 37381 91366 37408
rect 40824 37325 46844 37381
rect 46900 37325 53172 37381
rect 53228 37325 59500 37381
rect 59556 37325 65828 37381
rect 65884 37325 72156 37381
rect 72212 37325 78484 37381
rect 78540 37325 84812 37381
rect 84868 37325 91140 37381
rect 91196 37325 91366 37381
rect 40824 37296 91366 37325
rect 91478 37296 91560 37408
rect 40824 37240 91560 37296
rect 91672 37128 92008 40488
rect 40824 36904 92008 37128
rect 41160 36827 41272 36848
rect 41160 36771 41187 36827
rect 41243 36771 41272 36827
rect 41160 35560 41272 36771
rect 41328 36825 41440 36848
rect 41328 36769 41361 36825
rect 41417 36769 41440 36825
rect 41328 36396 41440 36769
rect 41328 36320 41709 36396
rect 46348 36218 46424 36904
rect 46816 36821 46928 36848
rect 46816 36765 46844 36821
rect 46900 36765 46928 36821
rect 46816 36736 46928 36765
rect 47488 36822 47600 36848
rect 47488 36766 47514 36822
rect 47570 36766 47600 36822
rect 46830 36218 46906 36736
rect 47488 35560 47600 36766
rect 47656 36813 47768 36848
rect 47656 36757 47684 36813
rect 47740 36757 47768 36813
rect 47656 36396 47768 36757
rect 47656 36320 48037 36396
rect 52676 36218 52752 36904
rect 53144 36821 53256 36848
rect 53144 36765 53172 36821
rect 53228 36765 53256 36821
rect 53144 36736 53256 36765
rect 53816 36817 53928 36848
rect 53816 36761 53844 36817
rect 53900 36761 53928 36817
rect 53158 36218 53234 36736
rect 53816 35560 53928 36761
rect 53984 36824 54096 36848
rect 53984 36768 54016 36824
rect 54072 36768 54096 36824
rect 53984 36396 54096 36768
rect 53984 36320 54365 36396
rect 59004 36218 59080 36904
rect 59472 36821 59584 36848
rect 59472 36765 59500 36821
rect 59556 36765 59584 36821
rect 59472 36736 59584 36765
rect 60144 36816 60256 36848
rect 60144 36760 60174 36816
rect 60230 36760 60256 36816
rect 59486 36218 59562 36736
rect 60144 35560 60256 36760
rect 60312 36821 60424 36848
rect 60312 36765 60339 36821
rect 60395 36765 60424 36821
rect 60312 36396 60424 36765
rect 60312 36320 60693 36396
rect 65332 36218 65408 36904
rect 65800 36821 65912 36848
rect 65800 36765 65828 36821
rect 65884 36765 65912 36821
rect 65800 36736 65912 36765
rect 66472 36823 66584 36848
rect 66472 36767 66499 36823
rect 66555 36767 66584 36823
rect 65814 36218 65890 36736
rect 66472 35560 66584 36767
rect 66640 36820 66752 36848
rect 66640 36764 66668 36820
rect 66724 36764 66752 36820
rect 66640 36396 66752 36764
rect 66640 36320 67021 36396
rect 71660 36218 71736 36904
rect 72128 36821 72240 36848
rect 72128 36765 72156 36821
rect 72212 36765 72240 36821
rect 72128 36736 72240 36765
rect 72800 36820 72912 36848
rect 72800 36764 72827 36820
rect 72883 36764 72912 36820
rect 72142 36218 72218 36736
rect 72800 35560 72912 36764
rect 72968 36816 73080 36848
rect 72968 36760 72997 36816
rect 73053 36760 73080 36816
rect 72968 36396 73080 36760
rect 72968 36320 73349 36396
rect 77988 36218 78064 36904
rect 78456 36821 78568 36848
rect 78456 36765 78484 36821
rect 78540 36765 78568 36821
rect 78456 36736 78568 36765
rect 79128 36817 79240 36848
rect 79128 36761 79155 36817
rect 79211 36761 79240 36817
rect 78470 36218 78546 36736
rect 79128 35560 79240 36761
rect 79296 36819 79408 36848
rect 79296 36763 79319 36819
rect 79375 36763 79408 36819
rect 79296 36396 79408 36763
rect 79296 36320 79677 36396
rect 84316 36218 84392 36904
rect 84784 36821 84896 36848
rect 84784 36765 84812 36821
rect 84868 36765 84896 36821
rect 84784 36736 84896 36765
rect 85456 36819 85568 36848
rect 85456 36763 85482 36819
rect 85538 36763 85568 36819
rect 84798 36218 84874 36736
rect 85456 35560 85568 36763
rect 85624 36820 85736 36848
rect 85624 36764 85655 36820
rect 85711 36764 85736 36820
rect 85624 36396 85736 36764
rect 85624 36320 86005 36396
rect 90644 36218 90720 36904
rect 91112 36821 91224 36848
rect 91112 36765 91140 36821
rect 91196 36765 91224 36821
rect 91112 36736 91224 36765
rect 91126 36218 91202 36736
rect 41160 35448 41749 35560
rect 47488 35448 48077 35560
rect 53816 35448 54405 35560
rect 60144 35448 60733 35560
rect 66472 35448 67061 35560
rect 72800 35448 73389 35560
rect 79128 35448 79717 35560
rect 85456 35448 86045 35560
rect 40824 34832 91560 34888
rect 40824 34802 91360 34832
rect 40824 34746 46811 34802
rect 46867 34746 53139 34802
rect 53195 34746 59467 34802
rect 59523 34746 65795 34802
rect 65851 34746 72123 34802
rect 72179 34746 78451 34802
rect 78507 34746 84779 34802
rect 84835 34746 91107 34802
rect 91163 34746 91360 34802
rect 40824 34720 91360 34746
rect 91472 34720 91560 34832
rect 40824 34664 91560 34720
rect 40544 34496 91560 34552
rect 40544 34384 40631 34496
rect 40743 34472 91560 34496
rect 40743 34416 41188 34472
rect 41244 34469 47516 34472
rect 41244 34416 43429 34469
rect 40743 34413 43429 34416
rect 43485 34416 47516 34469
rect 47572 34469 53844 34472
rect 47572 34416 49757 34469
rect 43485 34413 49757 34416
rect 49813 34416 53844 34469
rect 53900 34469 60172 34472
rect 53900 34416 56085 34469
rect 49813 34413 56085 34416
rect 56141 34416 60172 34469
rect 60228 34469 66500 34472
rect 60228 34416 62413 34469
rect 56141 34413 62413 34416
rect 62469 34416 66500 34469
rect 66556 34469 72828 34472
rect 66556 34416 68741 34469
rect 62469 34413 68741 34416
rect 68797 34416 72828 34469
rect 72884 34469 79156 34472
rect 72884 34416 75069 34469
rect 68797 34413 75069 34416
rect 75125 34416 79156 34469
rect 79212 34469 85484 34472
rect 79212 34416 81397 34469
rect 75125 34413 81397 34416
rect 81453 34416 85484 34469
rect 85540 34469 91560 34472
rect 85540 34416 87725 34469
rect 81453 34413 87725 34416
rect 87781 34413 91560 34469
rect 40743 34384 91560 34413
rect 40544 34328 91560 34384
rect 40152 34132 91560 34216
rect 40152 34076 41357 34132
rect 41413 34076 47685 34132
rect 47741 34076 54013 34132
rect 54069 34076 60341 34132
rect 60397 34076 66669 34132
rect 66725 34076 72997 34132
rect 73053 34076 79325 34132
rect 79381 34076 85653 34132
rect 85709 34076 91560 34132
rect 40152 33992 91560 34076
rect 40152 30632 40488 33992
rect 40824 33824 91560 33880
rect 40824 33797 91359 33824
rect 40824 33741 46844 33797
rect 46900 33741 53172 33797
rect 53228 33741 59500 33797
rect 59556 33741 65828 33797
rect 65884 33741 72156 33797
rect 72212 33741 78484 33797
rect 78540 33741 84812 33797
rect 84868 33741 91140 33797
rect 91196 33741 91359 33797
rect 40824 33712 91359 33741
rect 91471 33712 91560 33824
rect 40824 33656 91560 33712
rect 91672 33544 92008 36904
rect 40824 33320 92008 33544
rect 41160 33240 41272 33264
rect 41160 33184 41190 33240
rect 41246 33184 41272 33240
rect 41160 31976 41272 33184
rect 41328 33234 41440 33264
rect 41328 33178 41361 33234
rect 41417 33178 41440 33234
rect 41328 32812 41440 33178
rect 41328 32736 41709 32812
rect 46348 32634 46424 33320
rect 46816 33237 46928 33264
rect 46816 33181 46844 33237
rect 46900 33181 46928 33237
rect 46816 33152 46928 33181
rect 47488 33233 47600 33264
rect 47488 33177 47516 33233
rect 47572 33177 47600 33233
rect 46830 32634 46906 33152
rect 47488 31976 47600 33177
rect 47656 33235 47768 33264
rect 47656 33179 47682 33235
rect 47738 33179 47768 33235
rect 47656 32812 47768 33179
rect 47656 32736 48037 32812
rect 52676 32634 52752 33320
rect 53144 33237 53256 33264
rect 53144 33181 53172 33237
rect 53228 33181 53256 33237
rect 53144 33152 53256 33181
rect 53816 33232 53928 33264
rect 53816 33176 53843 33232
rect 53899 33176 53928 33232
rect 53158 32634 53234 33152
rect 53816 31976 53928 33176
rect 53984 33235 54096 33264
rect 53984 33179 54014 33235
rect 54070 33179 54096 33235
rect 53984 32812 54096 33179
rect 53984 32736 54365 32812
rect 59004 32634 59080 33320
rect 59472 33237 59584 33264
rect 59472 33181 59500 33237
rect 59556 33181 59584 33237
rect 59472 33152 59584 33181
rect 60144 33237 60256 33264
rect 60144 33181 60173 33237
rect 60229 33181 60256 33237
rect 59486 32634 59562 33152
rect 60144 31976 60256 33181
rect 60312 33235 60424 33264
rect 60312 33179 60342 33235
rect 60398 33179 60424 33235
rect 60312 32812 60424 33179
rect 60312 32736 60693 32812
rect 65332 32634 65408 33320
rect 65800 33237 65912 33264
rect 65800 33181 65828 33237
rect 65884 33181 65912 33237
rect 65800 33152 65912 33181
rect 66472 33231 66584 33264
rect 66472 33175 66503 33231
rect 66559 33175 66584 33231
rect 65814 32634 65890 33152
rect 66472 31976 66584 33175
rect 66640 33233 66752 33264
rect 66640 33177 66668 33233
rect 66724 33177 66752 33233
rect 66640 32812 66752 33177
rect 66640 32736 67021 32812
rect 71660 32634 71736 33320
rect 72128 33237 72240 33264
rect 72128 33181 72156 33237
rect 72212 33181 72240 33237
rect 72128 33152 72240 33181
rect 72800 33234 72912 33264
rect 72800 33178 72829 33234
rect 72885 33178 72912 33234
rect 72142 32634 72218 33152
rect 72800 31976 72912 33178
rect 72968 33235 73080 33264
rect 72968 33179 73003 33235
rect 73059 33179 73080 33235
rect 72968 32812 73080 33179
rect 72968 32736 73349 32812
rect 77988 32634 78064 33320
rect 78456 33237 78568 33264
rect 78456 33181 78484 33237
rect 78540 33181 78568 33237
rect 78456 33152 78568 33181
rect 79128 33235 79240 33264
rect 79128 33179 79154 33235
rect 79210 33179 79240 33235
rect 78470 32634 78546 33152
rect 79128 31976 79240 33179
rect 79296 33231 79408 33264
rect 79296 33175 79331 33231
rect 79387 33175 79408 33231
rect 79296 32812 79408 33175
rect 79296 32736 79677 32812
rect 84316 32634 84392 33320
rect 84784 33237 84896 33264
rect 84784 33181 84812 33237
rect 84868 33181 84896 33237
rect 84784 33152 84896 33181
rect 85456 33233 85568 33264
rect 85456 33177 85479 33233
rect 85535 33177 85568 33233
rect 84798 32634 84874 33152
rect 85456 31976 85568 33177
rect 85624 33235 85736 33264
rect 85624 33179 85652 33235
rect 85708 33179 85736 33235
rect 85624 32812 85736 33179
rect 85624 32736 86005 32812
rect 90644 32634 90720 33320
rect 91112 33237 91224 33264
rect 91112 33181 91140 33237
rect 91196 33181 91224 33237
rect 91112 33152 91224 33181
rect 91126 32634 91202 33152
rect 41160 31864 41749 31976
rect 47488 31864 48077 31976
rect 53816 31864 54405 31976
rect 60144 31864 60733 31976
rect 66472 31864 67061 31976
rect 72800 31864 73389 31976
rect 79128 31864 79717 31976
rect 85456 31864 86045 31976
rect 40824 31248 91560 31304
rect 40824 31218 91362 31248
rect 40824 31162 46811 31218
rect 46867 31162 53139 31218
rect 53195 31162 59467 31218
rect 59523 31162 65795 31218
rect 65851 31162 72123 31218
rect 72179 31162 78451 31218
rect 78507 31162 84779 31218
rect 84835 31162 91107 31218
rect 91163 31162 91362 31218
rect 40824 31136 91362 31162
rect 91474 31136 91560 31248
rect 40824 31080 91560 31136
rect 40544 30912 91560 30968
rect 40544 30800 40628 30912
rect 40740 30888 91560 30912
rect 40740 30832 41188 30888
rect 41244 30885 47516 30888
rect 41244 30832 43429 30885
rect 40740 30829 43429 30832
rect 43485 30832 47516 30885
rect 47572 30885 53844 30888
rect 47572 30832 49757 30885
rect 43485 30829 49757 30832
rect 49813 30832 53844 30885
rect 53900 30885 60172 30888
rect 53900 30832 56085 30885
rect 49813 30829 56085 30832
rect 56141 30832 60172 30885
rect 60228 30885 66500 30888
rect 60228 30832 62413 30885
rect 56141 30829 62413 30832
rect 62469 30832 66500 30885
rect 66556 30885 72828 30888
rect 66556 30832 68741 30885
rect 62469 30829 68741 30832
rect 68797 30832 72828 30885
rect 72884 30885 79156 30888
rect 72884 30832 75069 30885
rect 68797 30829 75069 30832
rect 75125 30832 79156 30885
rect 79212 30885 85484 30888
rect 79212 30832 81397 30885
rect 75125 30829 81397 30832
rect 81453 30832 85484 30885
rect 85540 30885 91560 30888
rect 85540 30832 87725 30885
rect 81453 30829 87725 30832
rect 87781 30829 91560 30885
rect 40740 30800 91560 30829
rect 40544 30744 91560 30800
rect 40152 30548 91560 30632
rect 40152 30492 41357 30548
rect 41413 30492 47685 30548
rect 47741 30492 54013 30548
rect 54069 30492 60341 30548
rect 60397 30492 66669 30548
rect 66725 30492 72997 30548
rect 73053 30492 79325 30548
rect 79381 30492 85653 30548
rect 85709 30492 91560 30548
rect 40152 30408 91560 30492
rect 40152 27048 40488 30408
rect 40824 30240 91560 30296
rect 40824 30213 91365 30240
rect 40824 30157 46844 30213
rect 46900 30157 53172 30213
rect 53228 30157 59500 30213
rect 59556 30157 65828 30213
rect 65884 30157 72156 30213
rect 72212 30157 78484 30213
rect 78540 30157 84812 30213
rect 84868 30157 91140 30213
rect 91196 30157 91365 30213
rect 40824 30128 91365 30157
rect 91477 30128 91560 30240
rect 40824 30072 91560 30128
rect 91672 29960 92008 33320
rect 40824 29736 92008 29960
rect 41160 29652 41272 29680
rect 41160 29596 41188 29652
rect 41244 29596 41272 29652
rect 41160 28392 41272 29596
rect 41328 29650 41440 29680
rect 41328 29594 41358 29650
rect 41414 29594 41440 29650
rect 41328 29228 41440 29594
rect 41328 29152 41709 29228
rect 46348 29050 46424 29736
rect 46816 29653 46928 29680
rect 46816 29597 46844 29653
rect 46900 29597 46928 29653
rect 46816 29568 46928 29597
rect 47488 29645 47600 29680
rect 47488 29589 47511 29645
rect 47567 29589 47600 29645
rect 46830 29050 46906 29568
rect 47488 28392 47600 29589
rect 47656 29646 47768 29680
rect 47656 29590 47686 29646
rect 47742 29590 47768 29646
rect 47656 29228 47768 29590
rect 47656 29152 48037 29228
rect 52676 29050 52752 29736
rect 53144 29653 53256 29680
rect 53144 29597 53172 29653
rect 53228 29597 53256 29653
rect 53144 29568 53256 29597
rect 53816 29648 53928 29680
rect 53816 29592 53838 29648
rect 53894 29592 53928 29648
rect 53158 29050 53234 29568
rect 53816 28392 53928 29592
rect 53984 29652 54096 29680
rect 53984 29596 54014 29652
rect 54070 29596 54096 29652
rect 53984 29228 54096 29596
rect 53984 29152 54365 29228
rect 59004 29050 59080 29736
rect 59472 29653 59584 29680
rect 59472 29597 59500 29653
rect 59556 29597 59584 29653
rect 59472 29568 59584 29597
rect 60144 29660 60256 29680
rect 60144 29604 60180 29660
rect 60236 29604 60256 29660
rect 59486 29050 59562 29568
rect 60144 28392 60256 29604
rect 60312 29659 60424 29680
rect 60312 29603 60343 29659
rect 60399 29603 60424 29659
rect 60312 29228 60424 29603
rect 60312 29152 60693 29228
rect 65332 29050 65408 29736
rect 65800 29653 65912 29680
rect 65800 29597 65828 29653
rect 65884 29597 65912 29653
rect 65800 29568 65912 29597
rect 66472 29648 66584 29680
rect 66472 29592 66496 29648
rect 66552 29592 66584 29648
rect 65814 29050 65890 29568
rect 66472 28392 66584 29592
rect 66640 29650 66752 29680
rect 66640 29594 66666 29650
rect 66722 29594 66752 29650
rect 66640 29228 66752 29594
rect 66640 29152 67021 29228
rect 71660 29050 71736 29736
rect 72128 29653 72240 29680
rect 72128 29597 72156 29653
rect 72212 29597 72240 29653
rect 72128 29568 72240 29597
rect 72800 29650 72912 29680
rect 72800 29594 72824 29650
rect 72880 29594 72912 29650
rect 72142 29050 72218 29568
rect 72800 28392 72912 29594
rect 72968 29651 73080 29680
rect 72968 29595 72995 29651
rect 73051 29595 73080 29651
rect 72968 29228 73080 29595
rect 72968 29152 73349 29228
rect 77988 29050 78064 29736
rect 78456 29653 78568 29680
rect 78456 29597 78484 29653
rect 78540 29597 78568 29653
rect 78456 29568 78568 29597
rect 79128 29648 79240 29680
rect 79128 29592 79149 29648
rect 79205 29592 79240 29648
rect 78470 29050 78546 29568
rect 79128 28392 79240 29592
rect 79296 29652 79408 29680
rect 79296 29596 79323 29652
rect 79379 29596 79408 29652
rect 79296 29228 79408 29596
rect 79296 29152 79677 29228
rect 84316 29050 84392 29736
rect 84784 29653 84896 29680
rect 84784 29597 84812 29653
rect 84868 29597 84896 29653
rect 84784 29568 84896 29597
rect 85456 29652 85568 29680
rect 85456 29596 85483 29652
rect 85539 29596 85568 29652
rect 84798 29050 84874 29568
rect 85456 28392 85568 29596
rect 85624 29650 85736 29680
rect 85624 29594 85659 29650
rect 85715 29594 85736 29650
rect 85624 29228 85736 29594
rect 85624 29152 86005 29228
rect 90644 29050 90720 29736
rect 91112 29653 91224 29680
rect 91112 29597 91140 29653
rect 91196 29597 91224 29653
rect 91112 29568 91224 29597
rect 91126 29050 91202 29568
rect 41160 28280 41749 28392
rect 47488 28280 48077 28392
rect 53816 28280 54405 28392
rect 60144 28280 60733 28392
rect 66472 28280 67061 28392
rect 72800 28280 73389 28392
rect 79128 28280 79717 28392
rect 85456 28280 86045 28392
rect 40824 27664 91560 27720
rect 40824 27634 91364 27664
rect 40824 27578 46811 27634
rect 46867 27578 53139 27634
rect 53195 27578 59467 27634
rect 59523 27578 65795 27634
rect 65851 27578 72123 27634
rect 72179 27578 78451 27634
rect 78507 27578 84779 27634
rect 84835 27578 91107 27634
rect 91163 27578 91364 27634
rect 40824 27552 91364 27578
rect 91476 27552 91560 27664
rect 40824 27496 91560 27552
rect 40544 27328 91560 27384
rect 40544 27216 40627 27328
rect 40739 27304 91560 27328
rect 40739 27248 41188 27304
rect 41244 27301 47516 27304
rect 41244 27248 43429 27301
rect 40739 27245 43429 27248
rect 43485 27248 47516 27301
rect 47572 27301 53844 27304
rect 47572 27248 49757 27301
rect 43485 27245 49757 27248
rect 49813 27248 53844 27301
rect 53900 27301 60172 27304
rect 53900 27248 56085 27301
rect 49813 27245 56085 27248
rect 56141 27248 60172 27301
rect 60228 27301 66500 27304
rect 60228 27248 62413 27301
rect 56141 27245 62413 27248
rect 62469 27248 66500 27301
rect 66556 27301 72828 27304
rect 66556 27248 68741 27301
rect 62469 27245 68741 27248
rect 68797 27248 72828 27301
rect 72884 27301 79156 27304
rect 72884 27248 75069 27301
rect 68797 27245 75069 27248
rect 75125 27248 79156 27301
rect 79212 27301 85484 27304
rect 79212 27248 81397 27301
rect 75125 27245 81397 27248
rect 81453 27248 85484 27301
rect 85540 27301 91560 27304
rect 85540 27248 87725 27301
rect 81453 27245 87725 27248
rect 87781 27245 91560 27301
rect 40739 27216 91560 27245
rect 40544 27160 91560 27216
rect 40152 26964 91560 27048
rect 40152 26908 41357 26964
rect 41413 26908 47685 26964
rect 47741 26908 54013 26964
rect 54069 26908 60341 26964
rect 60397 26908 66669 26964
rect 66725 26908 72997 26964
rect 73053 26908 79325 26964
rect 79381 26908 85653 26964
rect 85709 26908 91560 26964
rect 40152 26824 91560 26908
rect 40152 23464 40488 26824
rect 40824 26656 91560 26712
rect 40824 26629 91364 26656
rect 40824 26573 46844 26629
rect 46900 26573 53172 26629
rect 53228 26573 59500 26629
rect 59556 26573 65828 26629
rect 65884 26573 72156 26629
rect 72212 26573 78484 26629
rect 78540 26573 84812 26629
rect 84868 26573 91140 26629
rect 91196 26573 91364 26629
rect 40824 26544 91364 26573
rect 91476 26544 91560 26656
rect 40824 26488 91560 26544
rect 91672 26376 92008 29736
rect 40824 26152 92008 26376
rect 41160 26063 41272 26096
rect 41160 26007 41182 26063
rect 41238 26007 41272 26063
rect 41160 24808 41272 26007
rect 41328 26069 41440 26096
rect 41328 26013 41355 26069
rect 41411 26013 41440 26069
rect 41328 25644 41440 26013
rect 41328 25568 41709 25644
rect 46348 25466 46424 26152
rect 46816 26069 46928 26096
rect 46816 26013 46844 26069
rect 46900 26013 46928 26069
rect 46816 25984 46928 26013
rect 47488 26063 47600 26096
rect 47488 26007 47517 26063
rect 47573 26007 47600 26063
rect 46830 25466 46906 25984
rect 47488 24808 47600 26007
rect 47656 26066 47768 26096
rect 47656 26010 47685 26066
rect 47741 26010 47768 26066
rect 47656 25644 47768 26010
rect 47656 25568 48037 25644
rect 52676 25466 52752 26152
rect 53144 26069 53256 26096
rect 53144 26013 53172 26069
rect 53228 26013 53256 26069
rect 53144 25984 53256 26013
rect 53816 26064 53928 26096
rect 53816 26008 53846 26064
rect 53902 26008 53928 26064
rect 53158 25466 53234 25984
rect 53816 24808 53928 26008
rect 53984 26067 54096 26096
rect 53984 26011 54013 26067
rect 54069 26011 54096 26067
rect 53984 25644 54096 26011
rect 53984 25568 54365 25644
rect 59004 25466 59080 26152
rect 59472 26069 59584 26096
rect 59472 26013 59500 26069
rect 59556 26013 59584 26069
rect 59472 25984 59584 26013
rect 60144 26065 60256 26096
rect 60144 26009 60175 26065
rect 60231 26009 60256 26065
rect 59486 25466 59562 25984
rect 60144 24808 60256 26009
rect 60312 26068 60424 26096
rect 60312 26012 60341 26068
rect 60397 26012 60424 26068
rect 60312 25644 60424 26012
rect 60312 25568 60693 25644
rect 65332 25466 65408 26152
rect 65800 26069 65912 26096
rect 65800 26013 65828 26069
rect 65884 26013 65912 26069
rect 65800 25984 65912 26013
rect 66472 26066 66584 26096
rect 66472 26010 66499 26066
rect 66555 26010 66584 26066
rect 65814 25466 65890 25984
rect 66472 24808 66584 26010
rect 66640 26071 66752 26096
rect 66640 26015 66670 26071
rect 66726 26015 66752 26071
rect 66640 25644 66752 26015
rect 66640 25568 67021 25644
rect 71660 25466 71736 26152
rect 72128 26069 72240 26096
rect 72128 26013 72156 26069
rect 72212 26013 72240 26069
rect 72128 25984 72240 26013
rect 72800 26068 72912 26096
rect 72800 26012 72829 26068
rect 72885 26012 72912 26068
rect 72142 25466 72218 25984
rect 72800 24808 72912 26012
rect 72968 26067 73080 26096
rect 72968 26011 72998 26067
rect 73054 26011 73080 26067
rect 72968 25644 73080 26011
rect 72968 25568 73349 25644
rect 77988 25466 78064 26152
rect 78456 26069 78568 26096
rect 78456 26013 78484 26069
rect 78540 26013 78568 26069
rect 78456 25984 78568 26013
rect 79128 26071 79240 26096
rect 79128 26015 79156 26071
rect 79212 26015 79240 26071
rect 78470 25466 78546 25984
rect 79128 24808 79240 26015
rect 79296 26066 79408 26096
rect 79296 26010 79325 26066
rect 79381 26010 79408 26066
rect 79296 25644 79408 26010
rect 79296 25568 79677 25644
rect 84316 25466 84392 26152
rect 84784 26069 84896 26096
rect 84784 26013 84812 26069
rect 84868 26013 84896 26069
rect 84784 25984 84896 26013
rect 85456 26071 85568 26096
rect 85456 26015 85486 26071
rect 85542 26015 85568 26071
rect 84798 25466 84874 25984
rect 85456 24808 85568 26015
rect 85624 26068 85736 26096
rect 85624 26012 85655 26068
rect 85711 26012 85736 26068
rect 85624 25644 85736 26012
rect 85624 25568 86005 25644
rect 90644 25466 90720 26152
rect 91112 26069 91224 26096
rect 91112 26013 91140 26069
rect 91196 26013 91224 26069
rect 91112 25984 91224 26013
rect 91126 25466 91202 25984
rect 41160 24696 41749 24808
rect 47488 24696 48077 24808
rect 53816 24696 54405 24808
rect 60144 24696 60733 24808
rect 66472 24696 67061 24808
rect 72800 24696 73389 24808
rect 79128 24696 79717 24808
rect 85456 24696 86045 24808
rect 40824 24080 91560 24136
rect 40824 24050 91365 24080
rect 40824 23994 46811 24050
rect 46867 23994 53139 24050
rect 53195 23994 59467 24050
rect 59523 23994 65795 24050
rect 65851 23994 72123 24050
rect 72179 23994 78451 24050
rect 78507 23994 84779 24050
rect 84835 23994 91107 24050
rect 91163 23994 91365 24050
rect 40824 23968 91365 23994
rect 91477 23968 91560 24080
rect 40824 23912 91560 23968
rect 40544 23744 91560 23800
rect 40544 23632 40623 23744
rect 40735 23720 91560 23744
rect 40735 23664 41188 23720
rect 41244 23717 47516 23720
rect 41244 23664 43429 23717
rect 40735 23661 43429 23664
rect 43485 23664 47516 23717
rect 47572 23717 53844 23720
rect 47572 23664 49757 23717
rect 43485 23661 49757 23664
rect 49813 23664 53844 23717
rect 53900 23717 60172 23720
rect 53900 23664 56085 23717
rect 49813 23661 56085 23664
rect 56141 23664 60172 23717
rect 60228 23717 66500 23720
rect 60228 23664 62413 23717
rect 56141 23661 62413 23664
rect 62469 23664 66500 23717
rect 66556 23717 72828 23720
rect 66556 23664 68741 23717
rect 62469 23661 68741 23664
rect 68797 23664 72828 23717
rect 72884 23717 79156 23720
rect 72884 23664 75069 23717
rect 68797 23661 75069 23664
rect 75125 23664 79156 23717
rect 79212 23717 85484 23720
rect 79212 23664 81397 23717
rect 75125 23661 81397 23664
rect 81453 23664 85484 23717
rect 85540 23717 91560 23720
rect 85540 23664 87725 23717
rect 81453 23661 87725 23664
rect 87781 23661 91560 23717
rect 40735 23632 91560 23661
rect 40544 23576 91560 23632
rect 40152 23380 91560 23464
rect 40152 23324 41357 23380
rect 41413 23324 47685 23380
rect 47741 23324 54013 23380
rect 54069 23324 60341 23380
rect 60397 23324 66669 23380
rect 66725 23324 72997 23380
rect 73053 23324 79325 23380
rect 79381 23324 85653 23380
rect 85709 23324 91560 23380
rect 40152 23240 91560 23324
rect 40152 19880 40488 23240
rect 40824 23072 91560 23128
rect 40824 23045 91363 23072
rect 40824 22989 46844 23045
rect 46900 22989 53172 23045
rect 53228 22989 59500 23045
rect 59556 22989 65828 23045
rect 65884 22989 72156 23045
rect 72212 22989 78484 23045
rect 78540 22989 84812 23045
rect 84868 22989 91140 23045
rect 91196 22989 91363 23045
rect 40824 22960 91363 22989
rect 91475 22960 91560 23072
rect 40824 22904 91560 22960
rect 91672 22792 92008 26152
rect 40824 22568 92008 22792
rect 41160 22486 41272 22512
rect 41160 22430 41184 22486
rect 41240 22430 41272 22486
rect 41160 21224 41272 22430
rect 41328 22492 41440 22512
rect 41328 22436 41352 22492
rect 41408 22436 41440 22492
rect 41328 22060 41440 22436
rect 41328 21984 41709 22060
rect 46348 21882 46424 22568
rect 46816 22485 46928 22512
rect 46816 22429 46844 22485
rect 46900 22429 46928 22485
rect 46816 22400 46928 22429
rect 47488 22484 47600 22512
rect 47488 22428 47516 22484
rect 47572 22428 47600 22484
rect 46830 21882 46906 22400
rect 47488 21224 47600 22428
rect 47656 22486 47768 22512
rect 47656 22430 47686 22486
rect 47742 22430 47768 22486
rect 47656 22060 47768 22430
rect 47656 21984 48037 22060
rect 52676 21882 52752 22568
rect 53144 22485 53256 22512
rect 53144 22429 53172 22485
rect 53228 22429 53256 22485
rect 53144 22400 53256 22429
rect 53816 22490 53928 22512
rect 53816 22434 53848 22490
rect 53904 22434 53928 22490
rect 53158 21882 53234 22400
rect 53816 21224 53928 22434
rect 53984 22486 54096 22512
rect 53984 22430 54016 22486
rect 54072 22430 54096 22486
rect 53984 22060 54096 22430
rect 53984 21984 54365 22060
rect 59004 21882 59080 22568
rect 59472 22485 59584 22512
rect 59472 22429 59500 22485
rect 59556 22429 59584 22485
rect 59472 22400 59584 22429
rect 60144 22479 60256 22512
rect 60144 22423 60164 22479
rect 60220 22423 60256 22479
rect 59486 21882 59562 22400
rect 60144 21224 60256 22423
rect 60312 22488 60424 22512
rect 60312 22432 60339 22488
rect 60395 22432 60424 22488
rect 60312 22060 60424 22432
rect 60312 21984 60693 22060
rect 65332 21882 65408 22568
rect 65800 22485 65912 22512
rect 65800 22429 65828 22485
rect 65884 22429 65912 22485
rect 65800 22400 65912 22429
rect 66472 22483 66584 22512
rect 66472 22427 66498 22483
rect 66554 22427 66584 22483
rect 65814 21882 65890 22400
rect 66472 21224 66584 22427
rect 66640 22488 66752 22512
rect 66640 22432 66666 22488
rect 66722 22432 66752 22488
rect 66640 22060 66752 22432
rect 66640 21984 67021 22060
rect 71660 21882 71736 22568
rect 72128 22485 72240 22512
rect 72128 22429 72156 22485
rect 72212 22429 72240 22485
rect 72128 22400 72240 22429
rect 72800 22487 72912 22512
rect 72800 22431 72832 22487
rect 72888 22431 72912 22487
rect 72142 21882 72218 22400
rect 72800 21224 72912 22431
rect 72968 22483 73080 22512
rect 72968 22427 72989 22483
rect 73045 22427 73080 22483
rect 72968 22060 73080 22427
rect 72968 21984 73349 22060
rect 77988 21882 78064 22568
rect 78456 22485 78568 22512
rect 78456 22429 78484 22485
rect 78540 22429 78568 22485
rect 78456 22400 78568 22429
rect 79128 22480 79240 22512
rect 79128 22424 79152 22480
rect 79208 22424 79240 22480
rect 78470 21882 78546 22400
rect 79128 21224 79240 22424
rect 79296 22483 79408 22512
rect 79296 22427 79323 22483
rect 79379 22427 79408 22483
rect 79296 22060 79408 22427
rect 79296 21984 79677 22060
rect 84316 21882 84392 22568
rect 84784 22485 84896 22512
rect 84784 22429 84812 22485
rect 84868 22429 84896 22485
rect 84784 22400 84896 22429
rect 85456 22480 85568 22512
rect 85456 22424 85481 22480
rect 85537 22424 85568 22480
rect 84798 21882 84874 22400
rect 85456 21224 85568 22424
rect 85624 22482 85736 22512
rect 85624 22426 85655 22482
rect 85711 22426 85736 22482
rect 85624 22060 85736 22426
rect 85624 21984 86005 22060
rect 90644 21882 90720 22568
rect 91112 22485 91224 22512
rect 91112 22429 91140 22485
rect 91196 22429 91224 22485
rect 91112 22400 91224 22429
rect 91126 21882 91202 22400
rect 41160 21112 41749 21224
rect 47488 21112 48077 21224
rect 53816 21112 54405 21224
rect 60144 21112 60733 21224
rect 66472 21112 67061 21224
rect 72800 21112 73389 21224
rect 79128 21112 79717 21224
rect 85456 21112 86045 21224
rect 40824 20496 91560 20552
rect 40824 20466 91363 20496
rect 40824 20410 46811 20466
rect 46867 20410 53139 20466
rect 53195 20410 59467 20466
rect 59523 20410 65795 20466
rect 65851 20410 72123 20466
rect 72179 20410 78451 20466
rect 78507 20410 84779 20466
rect 84835 20410 91107 20466
rect 91163 20410 91363 20466
rect 40824 20384 91363 20410
rect 91475 20384 91560 20496
rect 40824 20328 91560 20384
rect 40544 20160 91560 20216
rect 40544 20048 40630 20160
rect 40742 20136 91560 20160
rect 40742 20080 41188 20136
rect 41244 20133 47516 20136
rect 41244 20080 43429 20133
rect 40742 20077 43429 20080
rect 43485 20080 47516 20133
rect 47572 20133 53844 20136
rect 47572 20080 49757 20133
rect 43485 20077 49757 20080
rect 49813 20080 53844 20133
rect 53900 20133 60172 20136
rect 53900 20080 56085 20133
rect 49813 20077 56085 20080
rect 56141 20080 60172 20133
rect 60228 20133 66500 20136
rect 60228 20080 62413 20133
rect 56141 20077 62413 20080
rect 62469 20080 66500 20133
rect 66556 20133 72828 20136
rect 66556 20080 68741 20133
rect 62469 20077 68741 20080
rect 68797 20080 72828 20133
rect 72884 20133 79156 20136
rect 72884 20080 75069 20133
rect 68797 20077 75069 20080
rect 75125 20080 79156 20133
rect 79212 20133 85484 20136
rect 79212 20080 81397 20133
rect 75125 20077 81397 20080
rect 81453 20080 85484 20133
rect 85540 20133 91560 20136
rect 85540 20080 87725 20133
rect 81453 20077 87725 20080
rect 87781 20077 91560 20133
rect 40742 20048 91560 20077
rect 40544 19992 91560 20048
rect 40152 19796 91560 19880
rect 40152 19740 41357 19796
rect 41413 19740 47685 19796
rect 47741 19740 54013 19796
rect 54069 19740 60341 19796
rect 60397 19740 66669 19796
rect 66725 19740 72997 19796
rect 73053 19740 79325 19796
rect 79381 19740 85653 19796
rect 85709 19740 91560 19796
rect 40152 19656 91560 19740
rect 40152 16296 40488 19656
rect 40824 19488 91560 19544
rect 40824 19461 91365 19488
rect 40824 19405 46844 19461
rect 46900 19405 53172 19461
rect 53228 19405 59500 19461
rect 59556 19405 65828 19461
rect 65884 19405 72156 19461
rect 72212 19405 78484 19461
rect 78540 19405 84812 19461
rect 84868 19405 91140 19461
rect 91196 19405 91365 19461
rect 40824 19376 91365 19405
rect 91477 19376 91560 19488
rect 40824 19320 91560 19376
rect 91672 19208 92008 22568
rect 40824 18984 92008 19208
rect 41160 18898 41272 18928
rect 41160 18842 41186 18898
rect 41242 18842 41272 18898
rect 41160 17640 41272 18842
rect 41328 18898 41440 18928
rect 41328 18842 41350 18898
rect 41406 18842 41440 18898
rect 41328 18476 41440 18842
rect 41328 18400 41709 18476
rect 46348 18298 46424 18984
rect 46816 18901 46928 18928
rect 46816 18845 46844 18901
rect 46900 18845 46928 18901
rect 46816 18816 46928 18845
rect 47488 18899 47600 18928
rect 47488 18843 47515 18899
rect 47571 18843 47600 18899
rect 46830 18298 46906 18816
rect 47488 17640 47600 18843
rect 47656 18898 47768 18928
rect 47656 18842 47686 18898
rect 47742 18842 47768 18898
rect 47656 18476 47768 18842
rect 47656 18400 48037 18476
rect 52676 18298 52752 18984
rect 53144 18901 53256 18928
rect 53144 18845 53172 18901
rect 53228 18845 53256 18901
rect 53144 18816 53256 18845
rect 53816 18903 53928 18928
rect 53816 18847 53847 18903
rect 53903 18847 53928 18903
rect 53158 18298 53234 18816
rect 53816 17640 53928 18847
rect 53984 18899 54096 18928
rect 53984 18843 54010 18899
rect 54066 18843 54096 18899
rect 53984 18476 54096 18843
rect 53984 18400 54365 18476
rect 59004 18298 59080 18984
rect 59472 18901 59584 18928
rect 59472 18845 59500 18901
rect 59556 18845 59584 18901
rect 59472 18816 59584 18845
rect 60144 18898 60256 18928
rect 60144 18842 60174 18898
rect 60230 18842 60256 18898
rect 59486 18298 59562 18816
rect 60144 17640 60256 18842
rect 60312 18898 60424 18928
rect 60312 18842 60339 18898
rect 60395 18842 60424 18898
rect 60312 18476 60424 18842
rect 60312 18400 60693 18476
rect 65332 18298 65408 18984
rect 65800 18901 65912 18928
rect 65800 18845 65828 18901
rect 65884 18845 65912 18901
rect 65800 18816 65912 18845
rect 66472 18900 66584 18928
rect 66472 18844 66500 18900
rect 66556 18844 66584 18900
rect 65814 18298 65890 18816
rect 66472 17640 66584 18844
rect 66640 18899 66752 18928
rect 66640 18843 66667 18899
rect 66723 18843 66752 18899
rect 66640 18476 66752 18843
rect 66640 18400 67021 18476
rect 71660 18298 71736 18984
rect 72128 18901 72240 18928
rect 72128 18845 72156 18901
rect 72212 18845 72240 18901
rect 72128 18816 72240 18845
rect 72800 18899 72912 18928
rect 72800 18843 72830 18899
rect 72886 18843 72912 18899
rect 72142 18298 72218 18816
rect 72800 17640 72912 18843
rect 72968 18899 73080 18928
rect 72968 18843 72999 18899
rect 73055 18843 73080 18899
rect 72968 18476 73080 18843
rect 72968 18400 73349 18476
rect 77988 18298 78064 18984
rect 78456 18901 78568 18928
rect 78456 18845 78484 18901
rect 78540 18845 78568 18901
rect 78456 18816 78568 18845
rect 79128 18901 79240 18928
rect 79128 18845 79159 18901
rect 79215 18845 79240 18901
rect 78470 18298 78546 18816
rect 79128 17640 79240 18845
rect 79296 18900 79408 18928
rect 79296 18844 79327 18900
rect 79383 18844 79408 18900
rect 79296 18476 79408 18844
rect 79296 18400 79677 18476
rect 84316 18298 84392 18984
rect 84784 18901 84896 18928
rect 84784 18845 84812 18901
rect 84868 18845 84896 18901
rect 84784 18816 84896 18845
rect 85456 18904 85568 18928
rect 85456 18848 85487 18904
rect 85543 18848 85568 18904
rect 84798 18298 84874 18816
rect 85456 17640 85568 18848
rect 85624 18899 85736 18928
rect 85624 18843 85651 18899
rect 85707 18843 85736 18899
rect 85624 18476 85736 18843
rect 85624 18400 86005 18476
rect 90644 18298 90720 18984
rect 91112 18901 91224 18928
rect 91112 18845 91140 18901
rect 91196 18845 91224 18901
rect 91112 18816 91224 18845
rect 91126 18298 91202 18816
rect 41160 17528 41749 17640
rect 47488 17528 48077 17640
rect 53816 17528 54405 17640
rect 60144 17528 60733 17640
rect 66472 17528 67061 17640
rect 72800 17528 73389 17640
rect 79128 17528 79717 17640
rect 85456 17528 86045 17640
rect 40824 16912 91560 16968
rect 40824 16882 91362 16912
rect 40824 16826 46811 16882
rect 46867 16826 53139 16882
rect 53195 16826 59467 16882
rect 59523 16826 65795 16882
rect 65851 16826 72123 16882
rect 72179 16826 78451 16882
rect 78507 16826 84779 16882
rect 84835 16826 91107 16882
rect 91163 16826 91362 16882
rect 40824 16800 91362 16826
rect 91474 16800 91560 16912
rect 40824 16744 91560 16800
rect 40544 16576 91560 16632
rect 40544 16464 40626 16576
rect 40738 16552 91560 16576
rect 40738 16496 41188 16552
rect 41244 16549 47516 16552
rect 41244 16496 43429 16549
rect 40738 16493 43429 16496
rect 43485 16496 47516 16549
rect 47572 16549 53844 16552
rect 47572 16496 49757 16549
rect 43485 16493 49757 16496
rect 49813 16496 53844 16549
rect 53900 16549 60172 16552
rect 53900 16496 56085 16549
rect 49813 16493 56085 16496
rect 56141 16496 60172 16549
rect 60228 16549 66500 16552
rect 60228 16496 62413 16549
rect 56141 16493 62413 16496
rect 62469 16496 66500 16549
rect 66556 16549 72828 16552
rect 66556 16496 68741 16549
rect 62469 16493 68741 16496
rect 68797 16496 72828 16549
rect 72884 16549 79156 16552
rect 72884 16496 75069 16549
rect 68797 16493 75069 16496
rect 75125 16496 79156 16549
rect 79212 16549 85484 16552
rect 79212 16496 81397 16549
rect 75125 16493 81397 16496
rect 81453 16496 85484 16549
rect 85540 16549 91560 16552
rect 85540 16496 87725 16549
rect 81453 16493 87725 16496
rect 87781 16493 91560 16549
rect 40738 16464 91560 16493
rect 40544 16408 91560 16464
rect 40152 16212 91560 16296
rect 40152 16156 41357 16212
rect 41413 16156 47685 16212
rect 47741 16156 54013 16212
rect 54069 16156 60341 16212
rect 60397 16156 66669 16212
rect 66725 16156 72997 16212
rect 73053 16156 79325 16212
rect 79381 16156 85653 16212
rect 85709 16156 91560 16212
rect 40152 16072 91560 16156
rect 40152 12712 40488 16072
rect 40824 15904 91560 15960
rect 40824 15877 91356 15904
rect 40824 15821 46844 15877
rect 46900 15821 53172 15877
rect 53228 15821 59500 15877
rect 59556 15821 65828 15877
rect 65884 15821 72156 15877
rect 72212 15821 78484 15877
rect 78540 15821 84812 15877
rect 84868 15821 91140 15877
rect 91196 15821 91356 15877
rect 40824 15792 91356 15821
rect 91468 15792 91560 15904
rect 40824 15736 91560 15792
rect 91672 15624 92008 18984
rect 40824 15400 92008 15624
rect 41160 15316 41272 15344
rect 41160 15260 41184 15316
rect 41240 15260 41272 15316
rect 41160 14056 41272 15260
rect 41328 15313 41440 15344
rect 41328 15257 41356 15313
rect 41412 15257 41440 15313
rect 41328 14892 41440 15257
rect 41328 14816 41709 14892
rect 46348 14714 46424 15400
rect 46816 15317 46928 15344
rect 46816 15261 46844 15317
rect 46900 15261 46928 15317
rect 46816 15232 46928 15261
rect 47488 15314 47600 15344
rect 47488 15258 47514 15314
rect 47570 15258 47600 15314
rect 46830 14714 46906 15232
rect 47488 14056 47600 15258
rect 47656 15316 47768 15344
rect 47656 15260 47683 15316
rect 47739 15260 47768 15316
rect 47656 14892 47768 15260
rect 47656 14816 48037 14892
rect 52676 14714 52752 15400
rect 53144 15317 53256 15344
rect 53144 15261 53172 15317
rect 53228 15261 53256 15317
rect 53144 15232 53256 15261
rect 53816 15314 53928 15344
rect 53816 15258 53842 15314
rect 53898 15258 53928 15314
rect 53158 14714 53234 15232
rect 53816 14056 53928 15258
rect 53984 15316 54096 15344
rect 53984 15260 54013 15316
rect 54069 15260 54096 15316
rect 53984 14892 54096 15260
rect 53984 14816 54365 14892
rect 59004 14714 59080 15400
rect 59472 15317 59584 15344
rect 59472 15261 59500 15317
rect 59556 15261 59584 15317
rect 59472 15232 59584 15261
rect 60144 15309 60256 15344
rect 60144 15253 60166 15309
rect 60222 15253 60256 15309
rect 59486 14714 59562 15232
rect 60144 14056 60256 15253
rect 60312 15314 60424 15344
rect 60312 15258 60343 15314
rect 60399 15258 60424 15314
rect 60312 14892 60424 15258
rect 60312 14816 60693 14892
rect 65332 14714 65408 15400
rect 65800 15317 65912 15344
rect 65800 15261 65828 15317
rect 65884 15261 65912 15317
rect 65800 15232 65912 15261
rect 66472 15315 66584 15344
rect 66472 15259 66498 15315
rect 66554 15259 66584 15315
rect 65814 14714 65890 15232
rect 66472 14056 66584 15259
rect 66640 15316 66752 15344
rect 66640 15260 66665 15316
rect 66721 15260 66752 15316
rect 66640 14892 66752 15260
rect 66640 14816 67021 14892
rect 71660 14714 71736 15400
rect 72128 15317 72240 15344
rect 72128 15261 72156 15317
rect 72212 15261 72240 15317
rect 72128 15232 72240 15261
rect 72800 15318 72912 15344
rect 72800 15262 72829 15318
rect 72885 15262 72912 15318
rect 72142 14714 72218 15232
rect 72800 14056 72912 15262
rect 72968 15316 73080 15344
rect 72968 15260 72994 15316
rect 73050 15260 73080 15316
rect 72968 14892 73080 15260
rect 72968 14816 73349 14892
rect 77988 14714 78064 15400
rect 78456 15317 78568 15344
rect 78456 15261 78484 15317
rect 78540 15261 78568 15317
rect 78456 15232 78568 15261
rect 79128 15314 79240 15344
rect 79128 15258 79153 15314
rect 79209 15258 79240 15314
rect 78470 14714 78546 15232
rect 79128 14056 79240 15258
rect 79296 15313 79408 15344
rect 79296 15257 79325 15313
rect 79381 15257 79408 15313
rect 79296 14892 79408 15257
rect 79296 14816 79677 14892
rect 84316 14714 84392 15400
rect 84784 15317 84896 15344
rect 84784 15261 84812 15317
rect 84868 15261 84896 15317
rect 84784 15232 84896 15261
rect 85456 15310 85568 15344
rect 85456 15254 85479 15310
rect 85535 15254 85568 15310
rect 84798 14714 84874 15232
rect 85456 14056 85568 15254
rect 85624 15314 85736 15344
rect 85624 15258 85649 15314
rect 85705 15258 85736 15314
rect 85624 14892 85736 15258
rect 85624 14816 86005 14892
rect 90644 14714 90720 15400
rect 91112 15317 91224 15344
rect 91112 15261 91140 15317
rect 91196 15261 91224 15317
rect 91112 15232 91224 15261
rect 91126 14714 91202 15232
rect 41160 13944 41749 14056
rect 47488 13944 48077 14056
rect 53816 13944 54405 14056
rect 60144 13944 60733 14056
rect 66472 13944 67061 14056
rect 72800 13944 73389 14056
rect 79128 13944 79717 14056
rect 85456 13944 86045 14056
rect 40824 13328 91560 13384
rect 40824 13298 91366 13328
rect 40824 13242 46811 13298
rect 46867 13242 53139 13298
rect 53195 13242 59467 13298
rect 59523 13242 65795 13298
rect 65851 13242 72123 13298
rect 72179 13242 78451 13298
rect 78507 13242 84779 13298
rect 84835 13242 91107 13298
rect 91163 13242 91366 13298
rect 40824 13216 91366 13242
rect 91478 13216 91560 13328
rect 40824 13160 91560 13216
rect 40824 12992 91560 13048
rect 40824 12880 41746 12992
rect 41858 12880 43036 12992
rect 43148 12965 44497 12992
rect 43148 12909 43429 12965
rect 43485 12909 44497 12965
rect 43148 12880 44497 12909
rect 44609 12880 48071 12992
rect 48183 12880 49364 12992
rect 49476 12965 50820 12992
rect 49476 12909 49757 12965
rect 49813 12909 50820 12965
rect 49476 12880 50820 12909
rect 50932 12880 54399 12992
rect 54511 12880 55689 12992
rect 55801 12965 57144 12992
rect 55801 12909 56085 12965
rect 56141 12909 57144 12965
rect 55801 12880 57144 12909
rect 57256 12965 91560 12992
rect 57256 12909 62413 12965
rect 62469 12909 68741 12965
rect 68797 12909 75069 12965
rect 75125 12909 81397 12965
rect 81453 12909 87725 12965
rect 87781 12909 91560 12965
rect 57256 12880 91560 12909
rect 40824 12824 91560 12880
rect 91672 12768 92008 15400
rect 92120 40992 92456 42056
rect 92120 40880 92232 40992
rect 92344 40880 92456 40992
rect 92120 37408 92456 40880
rect 92120 37296 92232 37408
rect 92344 37296 92456 37408
rect 92120 33824 92456 37296
rect 92120 33712 92232 33824
rect 92344 33712 92456 33824
rect 92120 30240 92456 33712
rect 92120 30128 92232 30240
rect 92344 30128 92456 30240
rect 92120 26656 92456 30128
rect 92120 26544 92232 26656
rect 92344 26544 92456 26656
rect 92120 23072 92456 26544
rect 92120 22960 92232 23072
rect 92344 22960 92456 23072
rect 92120 19488 92456 22960
rect 92120 19376 92232 19488
rect 92344 19376 92456 19488
rect 92120 15904 92456 19376
rect 92120 15792 92232 15904
rect 92344 15792 92456 15904
rect 92120 12768 92456 15792
rect 92568 38416 92904 42056
rect 92568 38304 92680 38416
rect 92792 38304 92904 38416
rect 92568 34832 92904 38304
rect 92568 34720 92680 34832
rect 92792 34720 92904 34832
rect 92568 31248 92904 34720
rect 92568 31136 92680 31248
rect 92792 31136 92904 31248
rect 92568 27664 92904 31136
rect 92568 27552 92680 27664
rect 92792 27552 92904 27664
rect 92568 24080 92904 27552
rect 92568 23968 92680 24080
rect 92792 23968 92904 24080
rect 92568 20496 92904 23968
rect 92568 20384 92680 20496
rect 92792 20384 92904 20496
rect 92568 16912 92904 20384
rect 92568 16800 92680 16912
rect 92792 16800 92904 16912
rect 92568 13328 92904 16800
rect 92568 13216 92680 13328
rect 92792 13216 92904 13328
rect 92568 12768 92904 13216
<< via1 >>
rect 41188 41584 41244 41640
rect 42392 41552 42504 41664
rect 43756 41552 43868 41664
rect 45212 41552 45324 41664
rect 47516 41584 47572 41640
rect 48720 41552 48832 41664
rect 50088 41552 50200 41664
rect 51550 41552 51662 41664
rect 53844 41584 53900 41640
rect 55048 41552 55160 41664
rect 56416 41552 56528 41664
rect 57873 41552 57985 41664
rect 60172 41584 60228 41640
rect 61376 41552 61488 41664
rect 62746 41552 62858 41664
rect 64204 41552 64316 41664
rect 66500 41584 66556 41640
rect 67704 41552 67816 41664
rect 69077 41552 69189 41664
rect 70528 41552 70640 41664
rect 72828 41584 72884 41640
rect 74032 41552 74144 41664
rect 75403 41552 75515 41664
rect 76860 41552 76972 41664
rect 79156 41584 79212 41640
rect 80360 41552 80472 41664
rect 81734 41552 81846 41664
rect 83186 41552 83298 41664
rect 85231 41584 85288 41642
rect 41357 41244 41413 41300
rect 47685 41244 47741 41300
rect 54013 41244 54069 41300
rect 60341 41244 60397 41300
rect 66669 41244 66725 41300
rect 72997 41244 73053 41300
rect 79325 41244 79381 41300
rect 46844 40909 46900 40965
rect 53172 40909 53228 40965
rect 59500 40909 59556 40965
rect 65828 40909 65884 40965
rect 72156 40909 72212 40965
rect 78484 40909 78540 40965
rect 84812 40909 84868 40965
rect 91363 40880 91475 40992
rect 41189 40349 41245 40405
rect 41363 40349 41419 40405
rect 46844 40349 46900 40405
rect 47517 40344 47573 40400
rect 47685 40349 47741 40405
rect 53172 40349 53228 40405
rect 53841 40348 53897 40404
rect 54016 40349 54072 40405
rect 59500 40349 59556 40405
rect 60173 40350 60229 40406
rect 60344 40347 60400 40403
rect 65828 40349 65884 40405
rect 66501 40349 66557 40405
rect 66673 40349 66729 40405
rect 72156 40349 72212 40405
rect 72829 40349 72885 40405
rect 72997 40347 73053 40403
rect 78484 40349 78540 40405
rect 79158 40347 79214 40403
rect 79328 40344 79384 40400
rect 84812 40349 84868 40405
rect 43420 39009 43476 39065
rect 49748 39009 49804 39065
rect 56076 39009 56132 39065
rect 62404 39009 62460 39065
rect 68732 39009 68788 39065
rect 75060 39009 75116 39065
rect 81388 39009 81444 39065
rect 41926 38864 41982 38920
rect 48254 38864 48310 38920
rect 54582 38864 54638 38920
rect 60910 38864 60966 38920
rect 67238 38864 67294 38920
rect 73566 38864 73622 38920
rect 79894 38864 79950 38920
rect 46811 38330 46867 38386
rect 53139 38330 53195 38386
rect 59467 38330 59523 38386
rect 65795 38330 65851 38386
rect 72123 38330 72179 38386
rect 78451 38330 78507 38386
rect 84779 38330 84835 38386
rect 91363 38304 91475 38416
rect 40626 37968 40738 38080
rect 41188 38000 41244 38056
rect 43429 37997 43485 38053
rect 47516 38000 47572 38056
rect 49757 37997 49813 38053
rect 53844 38000 53900 38056
rect 56085 37997 56141 38053
rect 60172 38000 60228 38056
rect 62413 37997 62469 38053
rect 66500 38000 66556 38056
rect 68741 37997 68797 38053
rect 72828 38000 72884 38056
rect 75069 37997 75125 38053
rect 79156 38000 79212 38056
rect 81397 37997 81453 38053
rect 85484 38000 85540 38056
rect 41357 37660 41413 37716
rect 47685 37660 47741 37716
rect 54013 37660 54069 37716
rect 60341 37660 60397 37716
rect 66669 37660 66725 37716
rect 72997 37660 73053 37716
rect 79325 37660 79381 37716
rect 85653 37660 85709 37716
rect 46844 37325 46900 37381
rect 53172 37325 53228 37381
rect 59500 37325 59556 37381
rect 65828 37325 65884 37381
rect 72156 37325 72212 37381
rect 78484 37325 78540 37381
rect 84812 37325 84868 37381
rect 91140 37325 91196 37381
rect 91366 37296 91478 37408
rect 41187 36771 41243 36827
rect 41361 36769 41417 36825
rect 46844 36765 46900 36821
rect 47514 36766 47570 36822
rect 47684 36757 47740 36813
rect 53172 36765 53228 36821
rect 53844 36761 53900 36817
rect 54016 36768 54072 36824
rect 59500 36765 59556 36821
rect 60174 36760 60230 36816
rect 60339 36765 60395 36821
rect 65828 36765 65884 36821
rect 66499 36767 66555 36823
rect 66668 36764 66724 36820
rect 72156 36765 72212 36821
rect 72827 36764 72883 36820
rect 72997 36760 73053 36816
rect 78484 36765 78540 36821
rect 79155 36761 79211 36817
rect 79319 36763 79375 36819
rect 84812 36765 84868 36821
rect 85482 36763 85538 36819
rect 85655 36764 85711 36820
rect 91140 36765 91196 36821
rect 43420 35425 43476 35481
rect 49748 35425 49804 35481
rect 56076 35425 56132 35481
rect 62404 35425 62460 35481
rect 68732 35425 68788 35481
rect 75060 35425 75116 35481
rect 81388 35425 81444 35481
rect 87716 35425 87772 35481
rect 41926 35280 41982 35336
rect 48254 35280 48310 35336
rect 54582 35280 54638 35336
rect 60910 35280 60966 35336
rect 67238 35280 67294 35336
rect 73566 35280 73622 35336
rect 79894 35280 79950 35336
rect 86222 35280 86278 35336
rect 46811 34746 46867 34802
rect 53139 34746 53195 34802
rect 59467 34746 59523 34802
rect 65795 34746 65851 34802
rect 72123 34746 72179 34802
rect 78451 34746 78507 34802
rect 84779 34746 84835 34802
rect 91107 34746 91163 34802
rect 91360 34720 91472 34832
rect 40631 34384 40743 34496
rect 41188 34416 41244 34472
rect 43429 34413 43485 34469
rect 47516 34416 47572 34472
rect 49757 34413 49813 34469
rect 53844 34416 53900 34472
rect 56085 34413 56141 34469
rect 60172 34416 60228 34472
rect 62413 34413 62469 34469
rect 66500 34416 66556 34472
rect 68741 34413 68797 34469
rect 72828 34416 72884 34472
rect 75069 34413 75125 34469
rect 79156 34416 79212 34472
rect 81397 34413 81453 34469
rect 85484 34416 85540 34472
rect 87725 34413 87781 34469
rect 41357 34076 41413 34132
rect 47685 34076 47741 34132
rect 54013 34076 54069 34132
rect 60341 34076 60397 34132
rect 66669 34076 66725 34132
rect 72997 34076 73053 34132
rect 79325 34076 79381 34132
rect 85653 34076 85709 34132
rect 46844 33741 46900 33797
rect 53172 33741 53228 33797
rect 59500 33741 59556 33797
rect 65828 33741 65884 33797
rect 72156 33741 72212 33797
rect 78484 33741 78540 33797
rect 84812 33741 84868 33797
rect 91140 33741 91196 33797
rect 91359 33712 91471 33824
rect 41190 33184 41246 33240
rect 41361 33178 41417 33234
rect 46844 33181 46900 33237
rect 47516 33177 47572 33233
rect 47682 33179 47738 33235
rect 53172 33181 53228 33237
rect 53843 33176 53899 33232
rect 54014 33179 54070 33235
rect 59500 33181 59556 33237
rect 60173 33181 60229 33237
rect 60342 33179 60398 33235
rect 65828 33181 65884 33237
rect 66503 33175 66559 33231
rect 66668 33177 66724 33233
rect 72156 33181 72212 33237
rect 72829 33178 72885 33234
rect 73003 33179 73059 33235
rect 78484 33181 78540 33237
rect 79154 33179 79210 33235
rect 79331 33175 79387 33231
rect 84812 33181 84868 33237
rect 85479 33177 85535 33233
rect 85652 33179 85708 33235
rect 91140 33181 91196 33237
rect 43420 31841 43476 31897
rect 49748 31841 49804 31897
rect 56076 31841 56132 31897
rect 62404 31841 62460 31897
rect 68732 31841 68788 31897
rect 75060 31841 75116 31897
rect 81388 31841 81444 31897
rect 87716 31841 87772 31897
rect 41926 31696 41982 31752
rect 48254 31696 48310 31752
rect 54582 31696 54638 31752
rect 60910 31696 60966 31752
rect 67238 31696 67294 31752
rect 73566 31696 73622 31752
rect 79894 31696 79950 31752
rect 86222 31696 86278 31752
rect 46811 31162 46867 31218
rect 53139 31162 53195 31218
rect 59467 31162 59523 31218
rect 65795 31162 65851 31218
rect 72123 31162 72179 31218
rect 78451 31162 78507 31218
rect 84779 31162 84835 31218
rect 91107 31162 91163 31218
rect 91362 31136 91474 31248
rect 40628 30800 40740 30912
rect 41188 30832 41244 30888
rect 43429 30829 43485 30885
rect 47516 30832 47572 30888
rect 49757 30829 49813 30885
rect 53844 30832 53900 30888
rect 56085 30829 56141 30885
rect 60172 30832 60228 30888
rect 62413 30829 62469 30885
rect 66500 30832 66556 30888
rect 68741 30829 68797 30885
rect 72828 30832 72884 30888
rect 75069 30829 75125 30885
rect 79156 30832 79212 30888
rect 81397 30829 81453 30885
rect 85484 30832 85540 30888
rect 87725 30829 87781 30885
rect 41357 30492 41413 30548
rect 47685 30492 47741 30548
rect 54013 30492 54069 30548
rect 60341 30492 60397 30548
rect 66669 30492 66725 30548
rect 72997 30492 73053 30548
rect 79325 30492 79381 30548
rect 85653 30492 85709 30548
rect 46844 30157 46900 30213
rect 53172 30157 53228 30213
rect 59500 30157 59556 30213
rect 65828 30157 65884 30213
rect 72156 30157 72212 30213
rect 78484 30157 78540 30213
rect 84812 30157 84868 30213
rect 91140 30157 91196 30213
rect 91365 30128 91477 30240
rect 41188 29596 41244 29652
rect 41358 29594 41414 29650
rect 46844 29597 46900 29653
rect 47511 29589 47567 29645
rect 47686 29590 47742 29646
rect 53172 29597 53228 29653
rect 53838 29592 53894 29648
rect 54014 29596 54070 29652
rect 59500 29597 59556 29653
rect 60180 29604 60236 29660
rect 60343 29603 60399 29659
rect 65828 29597 65884 29653
rect 66496 29592 66552 29648
rect 66666 29594 66722 29650
rect 72156 29597 72212 29653
rect 72824 29594 72880 29650
rect 72995 29595 73051 29651
rect 78484 29597 78540 29653
rect 79149 29592 79205 29648
rect 79323 29596 79379 29652
rect 84812 29597 84868 29653
rect 85483 29596 85539 29652
rect 85659 29594 85715 29650
rect 91140 29597 91196 29653
rect 43420 28257 43476 28313
rect 49748 28257 49804 28313
rect 56076 28257 56132 28313
rect 62404 28257 62460 28313
rect 68732 28257 68788 28313
rect 75060 28257 75116 28313
rect 81388 28257 81444 28313
rect 87716 28257 87772 28313
rect 41926 28112 41982 28168
rect 48254 28112 48310 28168
rect 54582 28112 54638 28168
rect 60910 28112 60966 28168
rect 67238 28112 67294 28168
rect 73566 28112 73622 28168
rect 79894 28112 79950 28168
rect 86222 28112 86278 28168
rect 46811 27578 46867 27634
rect 53139 27578 53195 27634
rect 59467 27578 59523 27634
rect 65795 27578 65851 27634
rect 72123 27578 72179 27634
rect 78451 27578 78507 27634
rect 84779 27578 84835 27634
rect 91107 27578 91163 27634
rect 91364 27552 91476 27664
rect 40627 27216 40739 27328
rect 41188 27248 41244 27304
rect 43429 27245 43485 27301
rect 47516 27248 47572 27304
rect 49757 27245 49813 27301
rect 53844 27248 53900 27304
rect 56085 27245 56141 27301
rect 60172 27248 60228 27304
rect 62413 27245 62469 27301
rect 66500 27248 66556 27304
rect 68741 27245 68797 27301
rect 72828 27248 72884 27304
rect 75069 27245 75125 27301
rect 79156 27248 79212 27304
rect 81397 27245 81453 27301
rect 85484 27248 85540 27304
rect 87725 27245 87781 27301
rect 41357 26908 41413 26964
rect 47685 26908 47741 26964
rect 54013 26908 54069 26964
rect 60341 26908 60397 26964
rect 66669 26908 66725 26964
rect 72997 26908 73053 26964
rect 79325 26908 79381 26964
rect 85653 26908 85709 26964
rect 46844 26573 46900 26629
rect 53172 26573 53228 26629
rect 59500 26573 59556 26629
rect 65828 26573 65884 26629
rect 72156 26573 72212 26629
rect 78484 26573 78540 26629
rect 84812 26573 84868 26629
rect 91140 26573 91196 26629
rect 91364 26544 91476 26656
rect 41182 26007 41238 26063
rect 41355 26013 41411 26069
rect 46844 26013 46900 26069
rect 47517 26007 47573 26063
rect 47685 26010 47741 26066
rect 53172 26013 53228 26069
rect 53846 26008 53902 26064
rect 54013 26011 54069 26067
rect 59500 26013 59556 26069
rect 60175 26009 60231 26065
rect 60341 26012 60397 26068
rect 65828 26013 65884 26069
rect 66499 26010 66555 26066
rect 66670 26015 66726 26071
rect 72156 26013 72212 26069
rect 72829 26012 72885 26068
rect 72998 26011 73054 26067
rect 78484 26013 78540 26069
rect 79156 26015 79212 26071
rect 79325 26010 79381 26066
rect 84812 26013 84868 26069
rect 85486 26015 85542 26071
rect 85655 26012 85711 26068
rect 91140 26013 91196 26069
rect 43420 24673 43476 24729
rect 49748 24673 49804 24729
rect 56076 24673 56132 24729
rect 62404 24673 62460 24729
rect 68732 24673 68788 24729
rect 75060 24673 75116 24729
rect 81388 24673 81444 24729
rect 87716 24673 87772 24729
rect 41926 24528 41982 24584
rect 48254 24528 48310 24584
rect 54582 24528 54638 24584
rect 60910 24528 60966 24584
rect 67238 24528 67294 24584
rect 73566 24528 73622 24584
rect 79894 24528 79950 24584
rect 86222 24528 86278 24584
rect 46811 23994 46867 24050
rect 53139 23994 53195 24050
rect 59467 23994 59523 24050
rect 65795 23994 65851 24050
rect 72123 23994 72179 24050
rect 78451 23994 78507 24050
rect 84779 23994 84835 24050
rect 91107 23994 91163 24050
rect 91365 23968 91477 24080
rect 40623 23632 40735 23744
rect 41188 23664 41244 23720
rect 43429 23661 43485 23717
rect 47516 23664 47572 23720
rect 49757 23661 49813 23717
rect 53844 23664 53900 23720
rect 56085 23661 56141 23717
rect 60172 23664 60228 23720
rect 62413 23661 62469 23717
rect 66500 23664 66556 23720
rect 68741 23661 68797 23717
rect 72828 23664 72884 23720
rect 75069 23661 75125 23717
rect 79156 23664 79212 23720
rect 81397 23661 81453 23717
rect 85484 23664 85540 23720
rect 87725 23661 87781 23717
rect 41357 23324 41413 23380
rect 47685 23324 47741 23380
rect 54013 23324 54069 23380
rect 60341 23324 60397 23380
rect 66669 23324 66725 23380
rect 72997 23324 73053 23380
rect 79325 23324 79381 23380
rect 85653 23324 85709 23380
rect 46844 22989 46900 23045
rect 53172 22989 53228 23045
rect 59500 22989 59556 23045
rect 65828 22989 65884 23045
rect 72156 22989 72212 23045
rect 78484 22989 78540 23045
rect 84812 22989 84868 23045
rect 91140 22989 91196 23045
rect 91363 22960 91475 23072
rect 41184 22430 41240 22486
rect 41352 22436 41408 22492
rect 46844 22429 46900 22485
rect 47516 22428 47572 22484
rect 47686 22430 47742 22486
rect 53172 22429 53228 22485
rect 53848 22434 53904 22490
rect 54016 22430 54072 22486
rect 59500 22429 59556 22485
rect 60164 22423 60220 22479
rect 60339 22432 60395 22488
rect 65828 22429 65884 22485
rect 66498 22427 66554 22483
rect 66666 22432 66722 22488
rect 72156 22429 72212 22485
rect 72832 22431 72888 22487
rect 72989 22427 73045 22483
rect 78484 22429 78540 22485
rect 79152 22424 79208 22480
rect 79323 22427 79379 22483
rect 84812 22429 84868 22485
rect 85481 22424 85537 22480
rect 85655 22426 85711 22482
rect 91140 22429 91196 22485
rect 43420 21089 43476 21145
rect 49748 21089 49804 21145
rect 56076 21089 56132 21145
rect 62404 21089 62460 21145
rect 68732 21089 68788 21145
rect 75060 21089 75116 21145
rect 81388 21089 81444 21145
rect 87716 21089 87772 21145
rect 41926 20944 41982 21000
rect 48254 20944 48310 21000
rect 54582 20944 54638 21000
rect 60910 20944 60966 21000
rect 67238 20944 67294 21000
rect 73566 20944 73622 21000
rect 79894 20944 79950 21000
rect 86222 20944 86278 21000
rect 46811 20410 46867 20466
rect 53139 20410 53195 20466
rect 59467 20410 59523 20466
rect 65795 20410 65851 20466
rect 72123 20410 72179 20466
rect 78451 20410 78507 20466
rect 84779 20410 84835 20466
rect 91107 20410 91163 20466
rect 91363 20384 91475 20496
rect 40630 20048 40742 20160
rect 41188 20080 41244 20136
rect 43429 20077 43485 20133
rect 47516 20080 47572 20136
rect 49757 20077 49813 20133
rect 53844 20080 53900 20136
rect 56085 20077 56141 20133
rect 60172 20080 60228 20136
rect 62413 20077 62469 20133
rect 66500 20080 66556 20136
rect 68741 20077 68797 20133
rect 72828 20080 72884 20136
rect 75069 20077 75125 20133
rect 79156 20080 79212 20136
rect 81397 20077 81453 20133
rect 85484 20080 85540 20136
rect 87725 20077 87781 20133
rect 41357 19740 41413 19796
rect 47685 19740 47741 19796
rect 54013 19740 54069 19796
rect 60341 19740 60397 19796
rect 66669 19740 66725 19796
rect 72997 19740 73053 19796
rect 79325 19740 79381 19796
rect 85653 19740 85709 19796
rect 46844 19405 46900 19461
rect 53172 19405 53228 19461
rect 59500 19405 59556 19461
rect 65828 19405 65884 19461
rect 72156 19405 72212 19461
rect 78484 19405 78540 19461
rect 84812 19405 84868 19461
rect 91140 19405 91196 19461
rect 91365 19376 91477 19488
rect 41186 18842 41242 18898
rect 41350 18842 41406 18898
rect 46844 18845 46900 18901
rect 47515 18843 47571 18899
rect 47686 18842 47742 18898
rect 53172 18845 53228 18901
rect 53847 18847 53903 18903
rect 54010 18843 54066 18899
rect 59500 18845 59556 18901
rect 60174 18842 60230 18898
rect 60339 18842 60395 18898
rect 65828 18845 65884 18901
rect 66500 18844 66556 18900
rect 66667 18843 66723 18899
rect 72156 18845 72212 18901
rect 72830 18843 72886 18899
rect 72999 18843 73055 18899
rect 78484 18845 78540 18901
rect 79159 18845 79215 18901
rect 79327 18844 79383 18900
rect 84812 18845 84868 18901
rect 85487 18848 85543 18904
rect 85651 18843 85707 18899
rect 91140 18845 91196 18901
rect 43420 17505 43476 17561
rect 49748 17505 49804 17561
rect 56076 17505 56132 17561
rect 62404 17505 62460 17561
rect 68732 17505 68788 17561
rect 75060 17505 75116 17561
rect 81388 17505 81444 17561
rect 87716 17505 87772 17561
rect 41926 17360 41982 17416
rect 48254 17360 48310 17416
rect 54582 17360 54638 17416
rect 60910 17360 60966 17416
rect 67238 17360 67294 17416
rect 73566 17360 73622 17416
rect 79894 17360 79950 17416
rect 86222 17360 86278 17416
rect 46811 16826 46867 16882
rect 53139 16826 53195 16882
rect 59467 16826 59523 16882
rect 65795 16826 65851 16882
rect 72123 16826 72179 16882
rect 78451 16826 78507 16882
rect 84779 16826 84835 16882
rect 91107 16826 91163 16882
rect 91362 16800 91474 16912
rect 40626 16464 40738 16576
rect 41188 16496 41244 16552
rect 43429 16493 43485 16549
rect 47516 16496 47572 16552
rect 49757 16493 49813 16549
rect 53844 16496 53900 16552
rect 56085 16493 56141 16549
rect 60172 16496 60228 16552
rect 62413 16493 62469 16549
rect 66500 16496 66556 16552
rect 68741 16493 68797 16549
rect 72828 16496 72884 16552
rect 75069 16493 75125 16549
rect 79156 16496 79212 16552
rect 81397 16493 81453 16549
rect 85484 16496 85540 16552
rect 87725 16493 87781 16549
rect 41357 16156 41413 16212
rect 47685 16156 47741 16212
rect 54013 16156 54069 16212
rect 60341 16156 60397 16212
rect 66669 16156 66725 16212
rect 72997 16156 73053 16212
rect 79325 16156 79381 16212
rect 85653 16156 85709 16212
rect 46844 15821 46900 15877
rect 53172 15821 53228 15877
rect 59500 15821 59556 15877
rect 65828 15821 65884 15877
rect 72156 15821 72212 15877
rect 78484 15821 78540 15877
rect 84812 15821 84868 15877
rect 91140 15821 91196 15877
rect 91356 15792 91468 15904
rect 41184 15260 41240 15316
rect 41356 15257 41412 15313
rect 46844 15261 46900 15317
rect 47514 15258 47570 15314
rect 47683 15260 47739 15316
rect 53172 15261 53228 15317
rect 53842 15258 53898 15314
rect 54013 15260 54069 15316
rect 59500 15261 59556 15317
rect 60166 15253 60222 15309
rect 60343 15258 60399 15314
rect 65828 15261 65884 15317
rect 66498 15259 66554 15315
rect 66665 15260 66721 15316
rect 72156 15261 72212 15317
rect 72829 15262 72885 15318
rect 72994 15260 73050 15316
rect 78484 15261 78540 15317
rect 79153 15258 79209 15314
rect 79325 15257 79381 15313
rect 84812 15261 84868 15317
rect 85479 15254 85535 15310
rect 85649 15258 85705 15314
rect 91140 15261 91196 15317
rect 43420 13921 43476 13977
rect 49748 13921 49804 13977
rect 56076 13921 56132 13977
rect 62404 13921 62460 13977
rect 68732 13921 68788 13977
rect 75060 13921 75116 13977
rect 81388 13921 81444 13977
rect 87716 13921 87772 13977
rect 41926 13776 41982 13832
rect 48254 13776 48310 13832
rect 54582 13776 54638 13832
rect 60910 13776 60966 13832
rect 67238 13776 67294 13832
rect 73566 13776 73622 13832
rect 79894 13776 79950 13832
rect 86222 13776 86278 13832
rect 46811 13242 46867 13298
rect 53139 13242 53195 13298
rect 59467 13242 59523 13298
rect 65795 13242 65851 13298
rect 72123 13242 72179 13298
rect 78451 13242 78507 13298
rect 84779 13242 84835 13298
rect 91107 13242 91163 13298
rect 91366 13216 91478 13328
rect 41746 12880 41858 12992
rect 43036 12880 43148 12992
rect 43429 12909 43485 12965
rect 44497 12880 44609 12992
rect 48071 12880 48183 12992
rect 49364 12880 49476 12992
rect 49757 12909 49813 12965
rect 50820 12880 50932 12992
rect 54399 12880 54511 12992
rect 55689 12880 55801 12992
rect 56085 12909 56141 12965
rect 57144 12880 57256 12992
rect 62413 12909 62469 12965
rect 68741 12909 68797 12965
rect 75069 12909 75125 12965
rect 81397 12909 81453 12965
rect 87725 12909 87781 12965
rect 92232 40880 92344 40992
rect 92232 37296 92344 37408
rect 92232 33712 92344 33824
rect 92232 30128 92344 30240
rect 92232 26544 92344 26656
rect 92232 22960 92344 23072
rect 92232 19376 92344 19488
rect 92232 15792 92344 15904
rect 92680 38304 92792 38416
rect 92680 34720 92792 34832
rect 92680 31136 92792 31248
rect 92680 27552 92792 27664
rect 92680 23968 92792 24080
rect 92680 20384 92792 20496
rect 92680 16800 92792 16912
rect 92680 13216 92792 13328
<< metal2 >>
rect 40880 38976 41048 42000
rect 41160 41640 41272 41720
rect 41160 41584 41188 41640
rect 41244 41584 41272 41640
rect 41160 40405 41272 41584
rect 42279 41664 42623 41719
rect 42279 41552 42392 41664
rect 42504 41552 42623 41664
rect 42279 41495 42623 41552
rect 43649 41664 43993 41720
rect 43649 41552 43756 41664
rect 43868 41552 43993 41664
rect 43649 41496 43993 41552
rect 45104 41664 45448 41720
rect 45104 41552 45212 41664
rect 45324 41552 45448 41664
rect 45104 41496 45448 41552
rect 41160 40349 41189 40405
rect 41245 40349 41272 40405
rect 41160 40320 41272 40349
rect 41328 41300 41440 41384
rect 41328 41244 41357 41300
rect 41413 41244 41440 41300
rect 41328 40405 41440 41244
rect 41328 40349 41363 40405
rect 41419 40349 41440 40405
rect 41328 40320 41440 40349
rect 46816 40965 46928 41048
rect 46816 40909 46844 40965
rect 46900 40909 46928 40965
rect 46816 40405 46928 40909
rect 46816 40349 46844 40405
rect 46900 40349 46928 40405
rect 46816 40320 46928 40349
rect 43400 39065 43512 39070
rect 43400 39009 43420 39065
rect 43476 39009 43512 39065
rect 40880 38920 41992 38976
rect 40880 38864 41926 38920
rect 41982 38864 41992 38920
rect 40880 38808 41992 38864
rect 40544 38080 40824 38136
rect 40544 37968 40626 38080
rect 40738 37968 40824 38080
rect 40544 37912 40824 37968
rect 40880 35392 41048 38808
rect 41160 38056 41272 38136
rect 41160 38000 41188 38056
rect 41244 38000 41272 38056
rect 41160 36827 41272 38000
rect 43400 38053 43512 39009
rect 46797 38472 46873 39144
rect 47208 38976 47376 42000
rect 47488 41640 47600 41720
rect 47488 41584 47516 41640
rect 47572 41584 47600 41640
rect 47488 40400 47600 41584
rect 48607 41664 48951 41720
rect 48607 41552 48720 41664
rect 48832 41552 48951 41664
rect 48607 41496 48951 41552
rect 49977 41664 50321 41720
rect 49977 41552 50088 41664
rect 50200 41552 50321 41664
rect 49977 41496 50321 41552
rect 51432 41664 51776 41720
rect 51432 41552 51550 41664
rect 51662 41552 51776 41664
rect 51432 41496 51776 41552
rect 47488 40344 47517 40400
rect 47573 40344 47600 40400
rect 47488 40320 47600 40344
rect 47656 41300 47768 41384
rect 47656 41244 47685 41300
rect 47741 41244 47768 41300
rect 47656 40405 47768 41244
rect 47656 40349 47685 40405
rect 47741 40349 47768 40405
rect 47656 40320 47768 40349
rect 53144 40965 53256 41048
rect 53144 40909 53172 40965
rect 53228 40909 53256 40965
rect 53144 40405 53256 40909
rect 53144 40349 53172 40405
rect 53228 40349 53256 40405
rect 53144 40320 53256 40349
rect 49728 39065 49840 39070
rect 49728 39009 49748 39065
rect 49804 39009 49840 39065
rect 47208 38920 48320 38976
rect 47208 38864 48254 38920
rect 48310 38864 48320 38920
rect 47208 38808 48320 38864
rect 46780 38386 46892 38472
rect 46780 38330 46811 38386
rect 46867 38330 46892 38386
rect 46780 38248 46892 38330
rect 43400 37997 43429 38053
rect 43485 37997 43512 38053
rect 43400 37912 43512 37997
rect 41160 36771 41187 36827
rect 41243 36771 41272 36827
rect 41160 36736 41272 36771
rect 41328 37716 41440 37800
rect 41328 37660 41357 37716
rect 41413 37660 41440 37716
rect 41328 36825 41440 37660
rect 41328 36769 41361 36825
rect 41417 36769 41440 36825
rect 41328 36736 41440 36769
rect 46816 37381 46928 37464
rect 46816 37325 46844 37381
rect 46900 37325 46928 37381
rect 46816 36821 46928 37325
rect 46816 36765 46844 36821
rect 46900 36765 46928 36821
rect 46816 36736 46928 36765
rect 43400 35481 43512 35486
rect 43400 35425 43420 35481
rect 43476 35425 43512 35481
rect 40880 35336 41992 35392
rect 40880 35280 41926 35336
rect 41982 35280 41992 35336
rect 40880 35224 41992 35280
rect 40544 34496 40824 34552
rect 40544 34384 40631 34496
rect 40743 34384 40824 34496
rect 40544 34328 40824 34384
rect 40880 31808 41048 35224
rect 41160 34472 41272 34552
rect 41160 34416 41188 34472
rect 41244 34416 41272 34472
rect 41160 33240 41272 34416
rect 43400 34469 43512 35425
rect 46797 34888 46873 35560
rect 47208 35392 47376 38808
rect 47488 38056 47600 38136
rect 47488 38000 47516 38056
rect 47572 38000 47600 38056
rect 47488 36822 47600 38000
rect 49728 38053 49840 39009
rect 53125 38472 53201 39144
rect 53536 38976 53704 42000
rect 53816 41640 53928 41720
rect 53816 41584 53844 41640
rect 53900 41584 53928 41640
rect 53816 40404 53928 41584
rect 54935 41664 55279 41720
rect 54935 41552 55048 41664
rect 55160 41552 55279 41664
rect 54935 41496 55279 41552
rect 56305 41664 56649 41720
rect 56305 41552 56416 41664
rect 56528 41552 56649 41664
rect 56305 41496 56649 41552
rect 57760 41664 58104 41720
rect 57760 41552 57873 41664
rect 57985 41552 58104 41664
rect 57760 41496 58104 41552
rect 53816 40348 53841 40404
rect 53897 40348 53928 40404
rect 53816 40320 53928 40348
rect 53984 41300 54096 41384
rect 53984 41244 54013 41300
rect 54069 41244 54096 41300
rect 53984 40405 54096 41244
rect 53984 40349 54016 40405
rect 54072 40349 54096 40405
rect 53984 40320 54096 40349
rect 59472 40965 59584 41048
rect 59472 40909 59500 40965
rect 59556 40909 59584 40965
rect 59472 40405 59584 40909
rect 59472 40349 59500 40405
rect 59556 40349 59584 40405
rect 59472 40320 59584 40349
rect 56056 39065 56168 39070
rect 56056 39009 56076 39065
rect 56132 39009 56168 39065
rect 53536 38920 54648 38976
rect 53536 38864 54582 38920
rect 54638 38864 54648 38920
rect 53536 38808 54648 38864
rect 53108 38386 53220 38472
rect 53108 38330 53139 38386
rect 53195 38330 53220 38386
rect 53108 38248 53220 38330
rect 49728 37997 49757 38053
rect 49813 37997 49840 38053
rect 49728 37912 49840 37997
rect 47488 36766 47514 36822
rect 47570 36766 47600 36822
rect 47488 36736 47600 36766
rect 47656 37716 47768 37800
rect 47656 37660 47685 37716
rect 47741 37660 47768 37716
rect 47656 36813 47768 37660
rect 47656 36757 47684 36813
rect 47740 36757 47768 36813
rect 47656 36736 47768 36757
rect 53144 37381 53256 37464
rect 53144 37325 53172 37381
rect 53228 37325 53256 37381
rect 53144 36821 53256 37325
rect 53144 36765 53172 36821
rect 53228 36765 53256 36821
rect 53144 36736 53256 36765
rect 49728 35481 49840 35486
rect 49728 35425 49748 35481
rect 49804 35425 49840 35481
rect 47208 35336 48320 35392
rect 47208 35280 48254 35336
rect 48310 35280 48320 35336
rect 47208 35224 48320 35280
rect 46780 34802 46892 34888
rect 46780 34746 46811 34802
rect 46867 34746 46892 34802
rect 46780 34664 46892 34746
rect 43400 34413 43429 34469
rect 43485 34413 43512 34469
rect 43400 34328 43512 34413
rect 41160 33184 41190 33240
rect 41246 33184 41272 33240
rect 41160 33152 41272 33184
rect 41328 34132 41440 34216
rect 41328 34076 41357 34132
rect 41413 34076 41440 34132
rect 41328 33234 41440 34076
rect 41328 33178 41361 33234
rect 41417 33178 41440 33234
rect 41328 33152 41440 33178
rect 46816 33797 46928 33880
rect 46816 33741 46844 33797
rect 46900 33741 46928 33797
rect 46816 33237 46928 33741
rect 46816 33181 46844 33237
rect 46900 33181 46928 33237
rect 46816 33152 46928 33181
rect 43400 31897 43512 31902
rect 43400 31841 43420 31897
rect 43476 31841 43512 31897
rect 40880 31752 41992 31808
rect 40880 31696 41926 31752
rect 41982 31696 41992 31752
rect 40880 31640 41992 31696
rect 40544 30912 40824 30968
rect 40544 30800 40628 30912
rect 40740 30800 40824 30912
rect 40544 30744 40824 30800
rect 40880 28224 41048 31640
rect 41160 30888 41272 30968
rect 41160 30832 41188 30888
rect 41244 30832 41272 30888
rect 41160 29652 41272 30832
rect 43400 30885 43512 31841
rect 46797 31304 46873 31976
rect 47208 31808 47376 35224
rect 47488 34472 47600 34552
rect 47488 34416 47516 34472
rect 47572 34416 47600 34472
rect 47488 33233 47600 34416
rect 49728 34469 49840 35425
rect 53125 34888 53201 35560
rect 53536 35392 53704 38808
rect 53816 38056 53928 38136
rect 53816 38000 53844 38056
rect 53900 38000 53928 38056
rect 53816 36817 53928 38000
rect 56056 38053 56168 39009
rect 59453 38472 59529 39144
rect 59864 38976 60032 42000
rect 60144 41640 60256 41720
rect 60144 41584 60172 41640
rect 60228 41584 60256 41640
rect 60144 40406 60256 41584
rect 61263 41664 61607 41720
rect 61263 41552 61376 41664
rect 61488 41552 61607 41664
rect 61263 41496 61607 41552
rect 62633 41664 62977 41720
rect 62633 41552 62746 41664
rect 62858 41552 62977 41664
rect 62633 41496 62977 41552
rect 64088 41664 64432 41720
rect 64088 41552 64204 41664
rect 64316 41552 64432 41664
rect 64088 41496 64432 41552
rect 60144 40350 60173 40406
rect 60229 40350 60256 40406
rect 60144 40320 60256 40350
rect 60312 41300 60424 41384
rect 60312 41244 60341 41300
rect 60397 41244 60424 41300
rect 60312 40403 60424 41244
rect 60312 40347 60344 40403
rect 60400 40347 60424 40403
rect 60312 40320 60424 40347
rect 65800 40965 65912 41048
rect 65800 40909 65828 40965
rect 65884 40909 65912 40965
rect 65800 40405 65912 40909
rect 65800 40349 65828 40405
rect 65884 40349 65912 40405
rect 65800 40320 65912 40349
rect 62384 39065 62496 39070
rect 62384 39009 62404 39065
rect 62460 39009 62496 39065
rect 59864 38920 60976 38976
rect 59864 38864 60910 38920
rect 60966 38864 60976 38920
rect 59864 38808 60976 38864
rect 59436 38386 59548 38472
rect 59436 38330 59467 38386
rect 59523 38330 59548 38386
rect 59436 38248 59548 38330
rect 56056 37997 56085 38053
rect 56141 37997 56168 38053
rect 56056 37912 56168 37997
rect 53816 36761 53844 36817
rect 53900 36761 53928 36817
rect 53816 36736 53928 36761
rect 53984 37716 54096 37800
rect 53984 37660 54013 37716
rect 54069 37660 54096 37716
rect 53984 36824 54096 37660
rect 53984 36768 54016 36824
rect 54072 36768 54096 36824
rect 53984 36736 54096 36768
rect 59472 37381 59584 37464
rect 59472 37325 59500 37381
rect 59556 37325 59584 37381
rect 59472 36821 59584 37325
rect 59472 36765 59500 36821
rect 59556 36765 59584 36821
rect 59472 36736 59584 36765
rect 56056 35481 56168 35486
rect 56056 35425 56076 35481
rect 56132 35425 56168 35481
rect 53536 35336 54648 35392
rect 53536 35280 54582 35336
rect 54638 35280 54648 35336
rect 53536 35224 54648 35280
rect 53108 34802 53220 34888
rect 53108 34746 53139 34802
rect 53195 34746 53220 34802
rect 53108 34664 53220 34746
rect 49728 34413 49757 34469
rect 49813 34413 49840 34469
rect 49728 34328 49840 34413
rect 47488 33177 47516 33233
rect 47572 33177 47600 33233
rect 47488 33152 47600 33177
rect 47656 34132 47768 34216
rect 47656 34076 47685 34132
rect 47741 34076 47768 34132
rect 47656 33235 47768 34076
rect 47656 33179 47682 33235
rect 47738 33179 47768 33235
rect 47656 33152 47768 33179
rect 53144 33797 53256 33880
rect 53144 33741 53172 33797
rect 53228 33741 53256 33797
rect 53144 33237 53256 33741
rect 53144 33181 53172 33237
rect 53228 33181 53256 33237
rect 53144 33152 53256 33181
rect 49728 31897 49840 31902
rect 49728 31841 49748 31897
rect 49804 31841 49840 31897
rect 47208 31752 48320 31808
rect 47208 31696 48254 31752
rect 48310 31696 48320 31752
rect 47208 31640 48320 31696
rect 46780 31218 46892 31304
rect 46780 31162 46811 31218
rect 46867 31162 46892 31218
rect 46780 31080 46892 31162
rect 43400 30829 43429 30885
rect 43485 30829 43512 30885
rect 43400 30744 43512 30829
rect 41160 29596 41188 29652
rect 41244 29596 41272 29652
rect 41160 29568 41272 29596
rect 41328 30548 41440 30632
rect 41328 30492 41357 30548
rect 41413 30492 41440 30548
rect 41328 29650 41440 30492
rect 41328 29594 41358 29650
rect 41414 29594 41440 29650
rect 41328 29568 41440 29594
rect 46816 30213 46928 30296
rect 46816 30157 46844 30213
rect 46900 30157 46928 30213
rect 46816 29653 46928 30157
rect 46816 29597 46844 29653
rect 46900 29597 46928 29653
rect 46816 29568 46928 29597
rect 43400 28313 43512 28318
rect 43400 28257 43420 28313
rect 43476 28257 43512 28313
rect 40880 28168 41992 28224
rect 40880 28112 41926 28168
rect 41982 28112 41992 28168
rect 40880 28056 41992 28112
rect 40544 27328 40824 27384
rect 40544 27216 40627 27328
rect 40739 27216 40824 27328
rect 40544 27160 40824 27216
rect 40880 24640 41048 28056
rect 41160 27304 41272 27384
rect 41160 27248 41188 27304
rect 41244 27248 41272 27304
rect 41160 26063 41272 27248
rect 43400 27301 43512 28257
rect 46797 27720 46873 28392
rect 47208 28224 47376 31640
rect 47488 30888 47600 30968
rect 47488 30832 47516 30888
rect 47572 30832 47600 30888
rect 47488 29645 47600 30832
rect 49728 30885 49840 31841
rect 53125 31304 53201 31976
rect 53536 31808 53704 35224
rect 53816 34472 53928 34552
rect 53816 34416 53844 34472
rect 53900 34416 53928 34472
rect 53816 33232 53928 34416
rect 56056 34469 56168 35425
rect 59453 34888 59529 35560
rect 59864 35392 60032 38808
rect 60144 38056 60256 38136
rect 60144 38000 60172 38056
rect 60228 38000 60256 38056
rect 60144 36816 60256 38000
rect 62384 38053 62496 39009
rect 65781 38472 65857 39144
rect 66192 38976 66360 42000
rect 66472 41640 66584 41720
rect 66472 41584 66500 41640
rect 66556 41584 66584 41640
rect 66472 40405 66584 41584
rect 67591 41664 67935 41720
rect 67591 41552 67704 41664
rect 67816 41552 67935 41664
rect 67591 41496 67935 41552
rect 68961 41664 69305 41720
rect 68961 41552 69077 41664
rect 69189 41552 69305 41664
rect 68961 41496 69305 41552
rect 70416 41664 70760 41720
rect 70416 41552 70528 41664
rect 70640 41552 70760 41664
rect 70416 41496 70760 41552
rect 66472 40349 66501 40405
rect 66557 40349 66584 40405
rect 66472 40320 66584 40349
rect 66640 41300 66752 41384
rect 66640 41244 66669 41300
rect 66725 41244 66752 41300
rect 66640 40405 66752 41244
rect 66640 40349 66673 40405
rect 66729 40349 66752 40405
rect 66640 40320 66752 40349
rect 72128 40965 72240 41048
rect 72128 40909 72156 40965
rect 72212 40909 72240 40965
rect 72128 40405 72240 40909
rect 72128 40349 72156 40405
rect 72212 40349 72240 40405
rect 72128 40320 72240 40349
rect 68712 39065 68824 39070
rect 68712 39009 68732 39065
rect 68788 39009 68824 39065
rect 66192 38920 67304 38976
rect 66192 38864 67238 38920
rect 67294 38864 67304 38920
rect 66192 38808 67304 38864
rect 65764 38386 65876 38472
rect 65764 38330 65795 38386
rect 65851 38330 65876 38386
rect 65764 38248 65876 38330
rect 62384 37997 62413 38053
rect 62469 37997 62496 38053
rect 62384 37912 62496 37997
rect 60144 36760 60174 36816
rect 60230 36760 60256 36816
rect 60144 36736 60256 36760
rect 60312 37716 60424 37800
rect 60312 37660 60341 37716
rect 60397 37660 60424 37716
rect 60312 36821 60424 37660
rect 60312 36765 60339 36821
rect 60395 36765 60424 36821
rect 60312 36736 60424 36765
rect 65800 37381 65912 37464
rect 65800 37325 65828 37381
rect 65884 37325 65912 37381
rect 65800 36821 65912 37325
rect 65800 36765 65828 36821
rect 65884 36765 65912 36821
rect 65800 36736 65912 36765
rect 62384 35481 62496 35486
rect 62384 35425 62404 35481
rect 62460 35425 62496 35481
rect 59864 35336 60976 35392
rect 59864 35280 60910 35336
rect 60966 35280 60976 35336
rect 59864 35224 60976 35280
rect 59436 34802 59548 34888
rect 59436 34746 59467 34802
rect 59523 34746 59548 34802
rect 59436 34664 59548 34746
rect 56056 34413 56085 34469
rect 56141 34413 56168 34469
rect 56056 34328 56168 34413
rect 53816 33176 53843 33232
rect 53899 33176 53928 33232
rect 53816 33152 53928 33176
rect 53984 34132 54096 34216
rect 53984 34076 54013 34132
rect 54069 34076 54096 34132
rect 53984 33235 54096 34076
rect 53984 33179 54014 33235
rect 54070 33179 54096 33235
rect 53984 33152 54096 33179
rect 59472 33797 59584 33880
rect 59472 33741 59500 33797
rect 59556 33741 59584 33797
rect 59472 33237 59584 33741
rect 59472 33181 59500 33237
rect 59556 33181 59584 33237
rect 59472 33152 59584 33181
rect 56056 31897 56168 31902
rect 56056 31841 56076 31897
rect 56132 31841 56168 31897
rect 53536 31752 54648 31808
rect 53536 31696 54582 31752
rect 54638 31696 54648 31752
rect 53536 31640 54648 31696
rect 53108 31218 53220 31304
rect 53108 31162 53139 31218
rect 53195 31162 53220 31218
rect 53108 31080 53220 31162
rect 49728 30829 49757 30885
rect 49813 30829 49840 30885
rect 49728 30744 49840 30829
rect 47488 29589 47511 29645
rect 47567 29589 47600 29645
rect 47488 29568 47600 29589
rect 47656 30548 47768 30632
rect 47656 30492 47685 30548
rect 47741 30492 47768 30548
rect 47656 29646 47768 30492
rect 47656 29590 47686 29646
rect 47742 29590 47768 29646
rect 47656 29568 47768 29590
rect 53144 30213 53256 30296
rect 53144 30157 53172 30213
rect 53228 30157 53256 30213
rect 53144 29653 53256 30157
rect 53144 29597 53172 29653
rect 53228 29597 53256 29653
rect 53144 29568 53256 29597
rect 49728 28313 49840 28318
rect 49728 28257 49748 28313
rect 49804 28257 49840 28313
rect 47208 28168 48320 28224
rect 47208 28112 48254 28168
rect 48310 28112 48320 28168
rect 47208 28056 48320 28112
rect 46780 27634 46892 27720
rect 46780 27578 46811 27634
rect 46867 27578 46892 27634
rect 46780 27496 46892 27578
rect 43400 27245 43429 27301
rect 43485 27245 43512 27301
rect 43400 27160 43512 27245
rect 41160 26007 41182 26063
rect 41238 26007 41272 26063
rect 41160 25984 41272 26007
rect 41328 26964 41440 27048
rect 41328 26908 41357 26964
rect 41413 26908 41440 26964
rect 41328 26069 41440 26908
rect 41328 26013 41355 26069
rect 41411 26013 41440 26069
rect 41328 25984 41440 26013
rect 46816 26629 46928 26712
rect 46816 26573 46844 26629
rect 46900 26573 46928 26629
rect 46816 26069 46928 26573
rect 46816 26013 46844 26069
rect 46900 26013 46928 26069
rect 46816 25984 46928 26013
rect 43400 24729 43512 24734
rect 43400 24673 43420 24729
rect 43476 24673 43512 24729
rect 40880 24584 41992 24640
rect 40880 24528 41926 24584
rect 41982 24528 41992 24584
rect 40880 24472 41992 24528
rect 40544 23744 40824 23800
rect 40544 23632 40623 23744
rect 40735 23632 40824 23744
rect 40544 23576 40824 23632
rect 40880 21056 41048 24472
rect 41160 23720 41272 23800
rect 41160 23664 41188 23720
rect 41244 23664 41272 23720
rect 41160 22486 41272 23664
rect 43400 23717 43512 24673
rect 46797 24136 46873 24808
rect 47208 24640 47376 28056
rect 47488 27304 47600 27384
rect 47488 27248 47516 27304
rect 47572 27248 47600 27304
rect 47488 26063 47600 27248
rect 49728 27301 49840 28257
rect 53125 27720 53201 28392
rect 53536 28224 53704 31640
rect 53816 30888 53928 30968
rect 53816 30832 53844 30888
rect 53900 30832 53928 30888
rect 53816 29648 53928 30832
rect 56056 30885 56168 31841
rect 59453 31304 59529 31976
rect 59864 31808 60032 35224
rect 60144 34472 60256 34552
rect 60144 34416 60172 34472
rect 60228 34416 60256 34472
rect 60144 33237 60256 34416
rect 62384 34469 62496 35425
rect 65781 34888 65857 35560
rect 66192 35392 66360 38808
rect 66472 38056 66584 38136
rect 66472 38000 66500 38056
rect 66556 38000 66584 38056
rect 66472 36823 66584 38000
rect 68712 38053 68824 39009
rect 72109 38472 72185 39144
rect 72520 38976 72688 42000
rect 72800 41640 72912 41720
rect 72800 41584 72828 41640
rect 72884 41584 72912 41640
rect 72800 40405 72912 41584
rect 73919 41664 74263 41720
rect 73919 41552 74032 41664
rect 74144 41552 74263 41664
rect 73919 41496 74263 41552
rect 75289 41664 75633 41720
rect 75289 41552 75403 41664
rect 75515 41552 75633 41664
rect 75289 41496 75633 41552
rect 76744 41664 77088 41720
rect 76744 41552 76860 41664
rect 76972 41552 77088 41664
rect 76744 41496 77088 41552
rect 72800 40349 72829 40405
rect 72885 40349 72912 40405
rect 72800 40320 72912 40349
rect 72968 41300 73080 41384
rect 72968 41244 72997 41300
rect 73053 41244 73080 41300
rect 72968 40403 73080 41244
rect 72968 40347 72997 40403
rect 73053 40347 73080 40403
rect 72968 40320 73080 40347
rect 78456 40965 78568 41048
rect 78456 40909 78484 40965
rect 78540 40909 78568 40965
rect 78456 40405 78568 40909
rect 78456 40349 78484 40405
rect 78540 40349 78568 40405
rect 78456 40320 78568 40349
rect 75040 39065 75152 39070
rect 75040 39009 75060 39065
rect 75116 39009 75152 39065
rect 72520 38920 73632 38976
rect 72520 38864 73566 38920
rect 73622 38864 73632 38920
rect 72520 38808 73632 38864
rect 72092 38386 72204 38472
rect 72092 38330 72123 38386
rect 72179 38330 72204 38386
rect 72092 38248 72204 38330
rect 68712 37997 68741 38053
rect 68797 37997 68824 38053
rect 68712 37912 68824 37997
rect 66472 36767 66499 36823
rect 66555 36767 66584 36823
rect 66472 36736 66584 36767
rect 66640 37716 66752 37800
rect 66640 37660 66669 37716
rect 66725 37660 66752 37716
rect 66640 36820 66752 37660
rect 66640 36764 66668 36820
rect 66724 36764 66752 36820
rect 66640 36736 66752 36764
rect 72128 37381 72240 37464
rect 72128 37325 72156 37381
rect 72212 37325 72240 37381
rect 72128 36821 72240 37325
rect 72128 36765 72156 36821
rect 72212 36765 72240 36821
rect 72128 36736 72240 36765
rect 68712 35481 68824 35486
rect 68712 35425 68732 35481
rect 68788 35425 68824 35481
rect 66192 35336 67304 35392
rect 66192 35280 67238 35336
rect 67294 35280 67304 35336
rect 66192 35224 67304 35280
rect 65764 34802 65876 34888
rect 65764 34746 65795 34802
rect 65851 34746 65876 34802
rect 65764 34664 65876 34746
rect 62384 34413 62413 34469
rect 62469 34413 62496 34469
rect 62384 34328 62496 34413
rect 60144 33181 60173 33237
rect 60229 33181 60256 33237
rect 60144 33152 60256 33181
rect 60312 34132 60424 34216
rect 60312 34076 60341 34132
rect 60397 34076 60424 34132
rect 60312 33235 60424 34076
rect 60312 33179 60342 33235
rect 60398 33179 60424 33235
rect 60312 33152 60424 33179
rect 65800 33797 65912 33880
rect 65800 33741 65828 33797
rect 65884 33741 65912 33797
rect 65800 33237 65912 33741
rect 65800 33181 65828 33237
rect 65884 33181 65912 33237
rect 65800 33152 65912 33181
rect 62384 31897 62496 31902
rect 62384 31841 62404 31897
rect 62460 31841 62496 31897
rect 59864 31752 60976 31808
rect 59864 31696 60910 31752
rect 60966 31696 60976 31752
rect 59864 31640 60976 31696
rect 59436 31218 59548 31304
rect 59436 31162 59467 31218
rect 59523 31162 59548 31218
rect 59436 31080 59548 31162
rect 56056 30829 56085 30885
rect 56141 30829 56168 30885
rect 56056 30744 56168 30829
rect 53816 29592 53838 29648
rect 53894 29592 53928 29648
rect 53816 29568 53928 29592
rect 53984 30548 54096 30632
rect 53984 30492 54013 30548
rect 54069 30492 54096 30548
rect 53984 29652 54096 30492
rect 53984 29596 54014 29652
rect 54070 29596 54096 29652
rect 53984 29568 54096 29596
rect 59472 30213 59584 30296
rect 59472 30157 59500 30213
rect 59556 30157 59584 30213
rect 59472 29653 59584 30157
rect 59472 29597 59500 29653
rect 59556 29597 59584 29653
rect 59472 29568 59584 29597
rect 56056 28313 56168 28318
rect 56056 28257 56076 28313
rect 56132 28257 56168 28313
rect 53536 28168 54648 28224
rect 53536 28112 54582 28168
rect 54638 28112 54648 28168
rect 53536 28056 54648 28112
rect 53108 27634 53220 27720
rect 53108 27578 53139 27634
rect 53195 27578 53220 27634
rect 53108 27496 53220 27578
rect 49728 27245 49757 27301
rect 49813 27245 49840 27301
rect 49728 27160 49840 27245
rect 47488 26007 47517 26063
rect 47573 26007 47600 26063
rect 47488 25984 47600 26007
rect 47656 26964 47768 27048
rect 47656 26908 47685 26964
rect 47741 26908 47768 26964
rect 47656 26066 47768 26908
rect 47656 26010 47685 26066
rect 47741 26010 47768 26066
rect 47656 25984 47768 26010
rect 53144 26629 53256 26712
rect 53144 26573 53172 26629
rect 53228 26573 53256 26629
rect 53144 26069 53256 26573
rect 53144 26013 53172 26069
rect 53228 26013 53256 26069
rect 53144 25984 53256 26013
rect 49728 24729 49840 24734
rect 49728 24673 49748 24729
rect 49804 24673 49840 24729
rect 47208 24584 48320 24640
rect 47208 24528 48254 24584
rect 48310 24528 48320 24584
rect 47208 24472 48320 24528
rect 46780 24050 46892 24136
rect 46780 23994 46811 24050
rect 46867 23994 46892 24050
rect 46780 23912 46892 23994
rect 43400 23661 43429 23717
rect 43485 23661 43512 23717
rect 43400 23576 43512 23661
rect 41160 22430 41184 22486
rect 41240 22430 41272 22486
rect 41160 22400 41272 22430
rect 41328 23380 41440 23464
rect 41328 23324 41357 23380
rect 41413 23324 41440 23380
rect 41328 22492 41440 23324
rect 41328 22436 41352 22492
rect 41408 22436 41440 22492
rect 41328 22400 41440 22436
rect 46816 23045 46928 23128
rect 46816 22989 46844 23045
rect 46900 22989 46928 23045
rect 46816 22485 46928 22989
rect 46816 22429 46844 22485
rect 46900 22429 46928 22485
rect 46816 22400 46928 22429
rect 43400 21145 43512 21150
rect 43400 21089 43420 21145
rect 43476 21089 43512 21145
rect 40880 21000 41992 21056
rect 40880 20944 41926 21000
rect 41982 20944 41992 21000
rect 40880 20888 41992 20944
rect 40544 20160 40824 20216
rect 40544 20048 40630 20160
rect 40742 20048 40824 20160
rect 40544 19992 40824 20048
rect 40880 17472 41048 20888
rect 41160 20136 41272 20216
rect 41160 20080 41188 20136
rect 41244 20080 41272 20136
rect 41160 18898 41272 20080
rect 43400 20133 43512 21089
rect 46797 20552 46873 21224
rect 47208 21056 47376 24472
rect 47488 23720 47600 23800
rect 47488 23664 47516 23720
rect 47572 23664 47600 23720
rect 47488 22484 47600 23664
rect 49728 23717 49840 24673
rect 53125 24136 53201 24808
rect 53536 24640 53704 28056
rect 53816 27304 53928 27384
rect 53816 27248 53844 27304
rect 53900 27248 53928 27304
rect 53816 26064 53928 27248
rect 56056 27301 56168 28257
rect 59453 27720 59529 28392
rect 59864 28224 60032 31640
rect 60144 30888 60256 30968
rect 60144 30832 60172 30888
rect 60228 30832 60256 30888
rect 60144 29660 60256 30832
rect 62384 30885 62496 31841
rect 65781 31304 65857 31976
rect 66192 31808 66360 35224
rect 66472 34472 66584 34552
rect 66472 34416 66500 34472
rect 66556 34416 66584 34472
rect 66472 33231 66584 34416
rect 68712 34469 68824 35425
rect 72109 34888 72185 35560
rect 72520 35392 72688 38808
rect 72800 38056 72912 38136
rect 72800 38000 72828 38056
rect 72884 38000 72912 38056
rect 72800 36820 72912 38000
rect 75040 38053 75152 39009
rect 78437 38472 78513 39144
rect 78848 38976 79016 42000
rect 79128 41640 79240 41720
rect 79128 41584 79156 41640
rect 79212 41584 79240 41640
rect 79128 40403 79240 41584
rect 80247 41664 80591 41720
rect 80247 41552 80360 41664
rect 80472 41552 80591 41664
rect 80247 41496 80591 41552
rect 81617 41664 81961 41720
rect 81617 41552 81734 41664
rect 81846 41552 81961 41664
rect 81617 41496 81961 41552
rect 83072 41664 83416 41720
rect 83072 41552 83186 41664
rect 83298 41552 83416 41664
rect 83072 41496 83416 41552
rect 85176 41642 85344 41720
rect 85176 41584 85231 41642
rect 85288 41584 85344 41642
rect 79128 40347 79158 40403
rect 79214 40347 79240 40403
rect 79128 40320 79240 40347
rect 79296 41300 79408 41384
rect 79296 41244 79325 41300
rect 79381 41244 79408 41300
rect 79296 40400 79408 41244
rect 79296 40344 79328 40400
rect 79384 40344 79408 40400
rect 79296 40320 79408 40344
rect 84784 40965 84896 41048
rect 84784 40909 84812 40965
rect 84868 40909 84896 40965
rect 84784 40405 84896 40909
rect 84784 40349 84812 40405
rect 84868 40349 84896 40405
rect 84784 40320 84896 40349
rect 81368 39065 81480 39070
rect 81368 39009 81388 39065
rect 81444 39009 81480 39065
rect 78848 38920 79960 38976
rect 78848 38864 79894 38920
rect 79950 38864 79960 38920
rect 78848 38808 79960 38864
rect 78420 38386 78532 38472
rect 78420 38330 78451 38386
rect 78507 38330 78532 38386
rect 78420 38248 78532 38330
rect 75040 37997 75069 38053
rect 75125 37997 75152 38053
rect 75040 37912 75152 37997
rect 72800 36764 72827 36820
rect 72883 36764 72912 36820
rect 72800 36736 72912 36764
rect 72968 37716 73080 37800
rect 72968 37660 72997 37716
rect 73053 37660 73080 37716
rect 72968 36816 73080 37660
rect 72968 36760 72997 36816
rect 73053 36760 73080 36816
rect 72968 36736 73080 36760
rect 78456 37381 78568 37464
rect 78456 37325 78484 37381
rect 78540 37325 78568 37381
rect 78456 36821 78568 37325
rect 78456 36765 78484 36821
rect 78540 36765 78568 36821
rect 78456 36736 78568 36765
rect 75040 35481 75152 35486
rect 75040 35425 75060 35481
rect 75116 35425 75152 35481
rect 72520 35336 73632 35392
rect 72520 35280 73566 35336
rect 73622 35280 73632 35336
rect 72520 35224 73632 35280
rect 72092 34802 72204 34888
rect 72092 34746 72123 34802
rect 72179 34746 72204 34802
rect 72092 34664 72204 34746
rect 68712 34413 68741 34469
rect 68797 34413 68824 34469
rect 68712 34328 68824 34413
rect 66472 33175 66503 33231
rect 66559 33175 66584 33231
rect 66472 33152 66584 33175
rect 66640 34132 66752 34216
rect 66640 34076 66669 34132
rect 66725 34076 66752 34132
rect 66640 33233 66752 34076
rect 66640 33177 66668 33233
rect 66724 33177 66752 33233
rect 66640 33152 66752 33177
rect 72128 33797 72240 33880
rect 72128 33741 72156 33797
rect 72212 33741 72240 33797
rect 72128 33237 72240 33741
rect 72128 33181 72156 33237
rect 72212 33181 72240 33237
rect 72128 33152 72240 33181
rect 68712 31897 68824 31902
rect 68712 31841 68732 31897
rect 68788 31841 68824 31897
rect 66192 31752 67304 31808
rect 66192 31696 67238 31752
rect 67294 31696 67304 31752
rect 66192 31640 67304 31696
rect 65764 31218 65876 31304
rect 65764 31162 65795 31218
rect 65851 31162 65876 31218
rect 65764 31080 65876 31162
rect 62384 30829 62413 30885
rect 62469 30829 62496 30885
rect 62384 30744 62496 30829
rect 60144 29604 60180 29660
rect 60236 29604 60256 29660
rect 60144 29568 60256 29604
rect 60312 30548 60424 30632
rect 60312 30492 60341 30548
rect 60397 30492 60424 30548
rect 60312 29659 60424 30492
rect 60312 29603 60343 29659
rect 60399 29603 60424 29659
rect 60312 29568 60424 29603
rect 65800 30213 65912 30296
rect 65800 30157 65828 30213
rect 65884 30157 65912 30213
rect 65800 29653 65912 30157
rect 65800 29597 65828 29653
rect 65884 29597 65912 29653
rect 65800 29568 65912 29597
rect 62384 28313 62496 28318
rect 62384 28257 62404 28313
rect 62460 28257 62496 28313
rect 59864 28168 60976 28224
rect 59864 28112 60910 28168
rect 60966 28112 60976 28168
rect 59864 28056 60976 28112
rect 59436 27634 59548 27720
rect 59436 27578 59467 27634
rect 59523 27578 59548 27634
rect 59436 27496 59548 27578
rect 56056 27245 56085 27301
rect 56141 27245 56168 27301
rect 56056 27160 56168 27245
rect 53816 26008 53846 26064
rect 53902 26008 53928 26064
rect 53816 25984 53928 26008
rect 53984 26964 54096 27048
rect 53984 26908 54013 26964
rect 54069 26908 54096 26964
rect 53984 26067 54096 26908
rect 53984 26011 54013 26067
rect 54069 26011 54096 26067
rect 53984 25984 54096 26011
rect 59472 26629 59584 26712
rect 59472 26573 59500 26629
rect 59556 26573 59584 26629
rect 59472 26069 59584 26573
rect 59472 26013 59500 26069
rect 59556 26013 59584 26069
rect 59472 25984 59584 26013
rect 56056 24729 56168 24734
rect 56056 24673 56076 24729
rect 56132 24673 56168 24729
rect 53536 24584 54648 24640
rect 53536 24528 54582 24584
rect 54638 24528 54648 24584
rect 53536 24472 54648 24528
rect 53108 24050 53220 24136
rect 53108 23994 53139 24050
rect 53195 23994 53220 24050
rect 53108 23912 53220 23994
rect 49728 23661 49757 23717
rect 49813 23661 49840 23717
rect 49728 23576 49840 23661
rect 47488 22428 47516 22484
rect 47572 22428 47600 22484
rect 47488 22400 47600 22428
rect 47656 23380 47768 23464
rect 47656 23324 47685 23380
rect 47741 23324 47768 23380
rect 47656 22486 47768 23324
rect 47656 22430 47686 22486
rect 47742 22430 47768 22486
rect 47656 22400 47768 22430
rect 53144 23045 53256 23128
rect 53144 22989 53172 23045
rect 53228 22989 53256 23045
rect 53144 22485 53256 22989
rect 53144 22429 53172 22485
rect 53228 22429 53256 22485
rect 53144 22400 53256 22429
rect 49728 21145 49840 21150
rect 49728 21089 49748 21145
rect 49804 21089 49840 21145
rect 47208 21000 48320 21056
rect 47208 20944 48254 21000
rect 48310 20944 48320 21000
rect 47208 20888 48320 20944
rect 46780 20466 46892 20552
rect 46780 20410 46811 20466
rect 46867 20410 46892 20466
rect 46780 20328 46892 20410
rect 43400 20077 43429 20133
rect 43485 20077 43512 20133
rect 43400 19992 43512 20077
rect 41160 18842 41186 18898
rect 41242 18842 41272 18898
rect 41160 18816 41272 18842
rect 41328 19796 41440 19880
rect 41328 19740 41357 19796
rect 41413 19740 41440 19796
rect 41328 18898 41440 19740
rect 41328 18842 41350 18898
rect 41406 18842 41440 18898
rect 41328 18816 41440 18842
rect 46816 19461 46928 19544
rect 46816 19405 46844 19461
rect 46900 19405 46928 19461
rect 46816 18901 46928 19405
rect 46816 18845 46844 18901
rect 46900 18845 46928 18901
rect 46816 18816 46928 18845
rect 43400 17561 43512 17566
rect 43400 17505 43420 17561
rect 43476 17505 43512 17561
rect 40880 17416 41992 17472
rect 40880 17360 41926 17416
rect 41982 17360 41992 17416
rect 40880 17304 41992 17360
rect 40544 16576 40824 16632
rect 40544 16464 40626 16576
rect 40738 16464 40824 16576
rect 40544 16408 40824 16464
rect 40880 13888 41048 17304
rect 41160 16552 41272 16632
rect 41160 16496 41188 16552
rect 41244 16496 41272 16552
rect 41160 15316 41272 16496
rect 43400 16549 43512 17505
rect 46797 16968 46873 17640
rect 47208 17472 47376 20888
rect 47488 20136 47600 20216
rect 47488 20080 47516 20136
rect 47572 20080 47600 20136
rect 47488 18899 47600 20080
rect 49728 20133 49840 21089
rect 53125 20552 53201 21224
rect 53536 21056 53704 24472
rect 53816 23720 53928 23800
rect 53816 23664 53844 23720
rect 53900 23664 53928 23720
rect 53816 22490 53928 23664
rect 56056 23717 56168 24673
rect 59453 24136 59529 24808
rect 59864 24640 60032 28056
rect 60144 27304 60256 27384
rect 60144 27248 60172 27304
rect 60228 27248 60256 27304
rect 60144 26065 60256 27248
rect 62384 27301 62496 28257
rect 65781 27720 65857 28392
rect 66192 28224 66360 31640
rect 66472 30888 66584 30968
rect 66472 30832 66500 30888
rect 66556 30832 66584 30888
rect 66472 29648 66584 30832
rect 68712 30885 68824 31841
rect 72109 31304 72185 31976
rect 72520 31808 72688 35224
rect 72800 34472 72912 34552
rect 72800 34416 72828 34472
rect 72884 34416 72912 34472
rect 72800 33234 72912 34416
rect 75040 34469 75152 35425
rect 78437 34888 78513 35560
rect 78848 35392 79016 38808
rect 79128 38056 79240 38136
rect 79128 38000 79156 38056
rect 79212 38000 79240 38056
rect 79128 36817 79240 38000
rect 81368 38053 81480 39009
rect 84765 38472 84841 39144
rect 84748 38386 84860 38472
rect 84748 38330 84779 38386
rect 84835 38330 84860 38386
rect 84748 38248 84860 38330
rect 81368 37997 81397 38053
rect 81453 37997 81480 38053
rect 81368 37912 81480 37997
rect 79128 36761 79155 36817
rect 79211 36761 79240 36817
rect 79128 36736 79240 36761
rect 79296 37716 79408 37800
rect 79296 37660 79325 37716
rect 79381 37660 79408 37716
rect 79296 36819 79408 37660
rect 79296 36763 79319 36819
rect 79375 36763 79408 36819
rect 79296 36736 79408 36763
rect 84784 37381 84896 37464
rect 84784 37325 84812 37381
rect 84868 37325 84896 37381
rect 84784 36821 84896 37325
rect 84784 36765 84812 36821
rect 84868 36765 84896 36821
rect 84784 36736 84896 36765
rect 81368 35481 81480 35486
rect 81368 35425 81388 35481
rect 81444 35425 81480 35481
rect 78848 35336 79960 35392
rect 78848 35280 79894 35336
rect 79950 35280 79960 35336
rect 78848 35224 79960 35280
rect 78420 34802 78532 34888
rect 78420 34746 78451 34802
rect 78507 34746 78532 34802
rect 78420 34664 78532 34746
rect 75040 34413 75069 34469
rect 75125 34413 75152 34469
rect 75040 34328 75152 34413
rect 72800 33178 72829 33234
rect 72885 33178 72912 33234
rect 72800 33152 72912 33178
rect 72968 34132 73080 34216
rect 72968 34076 72997 34132
rect 73053 34076 73080 34132
rect 72968 33235 73080 34076
rect 72968 33179 73003 33235
rect 73059 33179 73080 33235
rect 72968 33152 73080 33179
rect 78456 33797 78568 33880
rect 78456 33741 78484 33797
rect 78540 33741 78568 33797
rect 78456 33237 78568 33741
rect 78456 33181 78484 33237
rect 78540 33181 78568 33237
rect 78456 33152 78568 33181
rect 75040 31897 75152 31902
rect 75040 31841 75060 31897
rect 75116 31841 75152 31897
rect 72520 31752 73632 31808
rect 72520 31696 73566 31752
rect 73622 31696 73632 31752
rect 72520 31640 73632 31696
rect 72092 31218 72204 31304
rect 72092 31162 72123 31218
rect 72179 31162 72204 31218
rect 72092 31080 72204 31162
rect 68712 30829 68741 30885
rect 68797 30829 68824 30885
rect 68712 30744 68824 30829
rect 66472 29592 66496 29648
rect 66552 29592 66584 29648
rect 66472 29568 66584 29592
rect 66640 30548 66752 30632
rect 66640 30492 66669 30548
rect 66725 30492 66752 30548
rect 66640 29650 66752 30492
rect 66640 29594 66666 29650
rect 66722 29594 66752 29650
rect 66640 29568 66752 29594
rect 72128 30213 72240 30296
rect 72128 30157 72156 30213
rect 72212 30157 72240 30213
rect 72128 29653 72240 30157
rect 72128 29597 72156 29653
rect 72212 29597 72240 29653
rect 72128 29568 72240 29597
rect 68712 28313 68824 28318
rect 68712 28257 68732 28313
rect 68788 28257 68824 28313
rect 66192 28168 67304 28224
rect 66192 28112 67238 28168
rect 67294 28112 67304 28168
rect 66192 28056 67304 28112
rect 65764 27634 65876 27720
rect 65764 27578 65795 27634
rect 65851 27578 65876 27634
rect 65764 27496 65876 27578
rect 62384 27245 62413 27301
rect 62469 27245 62496 27301
rect 62384 27160 62496 27245
rect 60144 26009 60175 26065
rect 60231 26009 60256 26065
rect 60144 25984 60256 26009
rect 60312 26964 60424 27048
rect 60312 26908 60341 26964
rect 60397 26908 60424 26964
rect 60312 26068 60424 26908
rect 60312 26012 60341 26068
rect 60397 26012 60424 26068
rect 60312 25984 60424 26012
rect 65800 26629 65912 26712
rect 65800 26573 65828 26629
rect 65884 26573 65912 26629
rect 65800 26069 65912 26573
rect 65800 26013 65828 26069
rect 65884 26013 65912 26069
rect 65800 25984 65912 26013
rect 62384 24729 62496 24734
rect 62384 24673 62404 24729
rect 62460 24673 62496 24729
rect 59864 24584 60976 24640
rect 59864 24528 60910 24584
rect 60966 24528 60976 24584
rect 59864 24472 60976 24528
rect 59436 24050 59548 24136
rect 59436 23994 59467 24050
rect 59523 23994 59548 24050
rect 59436 23912 59548 23994
rect 56056 23661 56085 23717
rect 56141 23661 56168 23717
rect 56056 23576 56168 23661
rect 53816 22434 53848 22490
rect 53904 22434 53928 22490
rect 53816 22400 53928 22434
rect 53984 23380 54096 23464
rect 53984 23324 54013 23380
rect 54069 23324 54096 23380
rect 53984 22486 54096 23324
rect 53984 22430 54016 22486
rect 54072 22430 54096 22486
rect 53984 22400 54096 22430
rect 59472 23045 59584 23128
rect 59472 22989 59500 23045
rect 59556 22989 59584 23045
rect 59472 22485 59584 22989
rect 59472 22429 59500 22485
rect 59556 22429 59584 22485
rect 59472 22400 59584 22429
rect 56056 21145 56168 21150
rect 56056 21089 56076 21145
rect 56132 21089 56168 21145
rect 53536 21000 54648 21056
rect 53536 20944 54582 21000
rect 54638 20944 54648 21000
rect 53536 20888 54648 20944
rect 53108 20466 53220 20552
rect 53108 20410 53139 20466
rect 53195 20410 53220 20466
rect 53108 20328 53220 20410
rect 49728 20077 49757 20133
rect 49813 20077 49840 20133
rect 49728 19992 49840 20077
rect 47488 18843 47515 18899
rect 47571 18843 47600 18899
rect 47488 18816 47600 18843
rect 47656 19796 47768 19880
rect 47656 19740 47685 19796
rect 47741 19740 47768 19796
rect 47656 18898 47768 19740
rect 47656 18842 47686 18898
rect 47742 18842 47768 18898
rect 47656 18816 47768 18842
rect 53144 19461 53256 19544
rect 53144 19405 53172 19461
rect 53228 19405 53256 19461
rect 53144 18901 53256 19405
rect 53144 18845 53172 18901
rect 53228 18845 53256 18901
rect 53144 18816 53256 18845
rect 49728 17561 49840 17566
rect 49728 17505 49748 17561
rect 49804 17505 49840 17561
rect 47208 17416 48320 17472
rect 47208 17360 48254 17416
rect 48310 17360 48320 17416
rect 47208 17304 48320 17360
rect 46780 16882 46892 16968
rect 46780 16826 46811 16882
rect 46867 16826 46892 16882
rect 46780 16744 46892 16826
rect 43400 16493 43429 16549
rect 43485 16493 43512 16549
rect 43400 16408 43512 16493
rect 41160 15260 41184 15316
rect 41240 15260 41272 15316
rect 41160 15232 41272 15260
rect 41328 16212 41440 16296
rect 41328 16156 41357 16212
rect 41413 16156 41440 16212
rect 41328 15313 41440 16156
rect 41328 15257 41356 15313
rect 41412 15257 41440 15313
rect 41328 15232 41440 15257
rect 46816 15877 46928 15960
rect 46816 15821 46844 15877
rect 46900 15821 46928 15877
rect 46816 15317 46928 15821
rect 46816 15261 46844 15317
rect 46900 15261 46928 15317
rect 46816 15232 46928 15261
rect 43400 13977 43512 13982
rect 43400 13921 43420 13977
rect 43476 13921 43512 13977
rect 40880 13832 41992 13888
rect 40880 13776 41926 13832
rect 41982 13776 41992 13832
rect 40880 13720 41992 13776
rect 40880 12656 41048 13720
rect 41630 12992 41974 13048
rect 41630 12880 41746 12992
rect 41858 12880 41974 12992
rect 41630 12824 41974 12880
rect 42922 12992 43266 13048
rect 42922 12880 43036 12992
rect 43148 12880 43266 12992
rect 42922 12824 43266 12880
rect 43400 12965 43512 13921
rect 46797 13384 46873 14056
rect 47208 13888 47376 17304
rect 47488 16552 47600 16632
rect 47488 16496 47516 16552
rect 47572 16496 47600 16552
rect 47488 15314 47600 16496
rect 49728 16549 49840 17505
rect 53125 16968 53201 17640
rect 53536 17472 53704 20888
rect 53816 20136 53928 20216
rect 53816 20080 53844 20136
rect 53900 20080 53928 20136
rect 53816 18903 53928 20080
rect 56056 20133 56168 21089
rect 59453 20552 59529 21224
rect 59864 21056 60032 24472
rect 60144 23720 60256 23800
rect 60144 23664 60172 23720
rect 60228 23664 60256 23720
rect 60144 22479 60256 23664
rect 62384 23717 62496 24673
rect 65781 24136 65857 24808
rect 66192 24640 66360 28056
rect 66472 27304 66584 27384
rect 66472 27248 66500 27304
rect 66556 27248 66584 27304
rect 66472 26066 66584 27248
rect 68712 27301 68824 28257
rect 72109 27720 72185 28392
rect 72520 28224 72688 31640
rect 72800 30888 72912 30968
rect 72800 30832 72828 30888
rect 72884 30832 72912 30888
rect 72800 29650 72912 30832
rect 75040 30885 75152 31841
rect 78437 31304 78513 31976
rect 78848 31808 79016 35224
rect 79128 34472 79240 34552
rect 79128 34416 79156 34472
rect 79212 34416 79240 34472
rect 79128 33235 79240 34416
rect 81368 34469 81480 35425
rect 84765 34888 84841 35560
rect 85176 35392 85344 41584
rect 91280 40992 92456 41048
rect 91280 40880 91363 40992
rect 91475 40880 92232 40992
rect 92344 40880 92456 40992
rect 91280 40824 92456 40880
rect 91280 38416 92904 38472
rect 91280 38304 91363 38416
rect 91475 38304 92680 38416
rect 92792 38304 92904 38416
rect 91280 38248 92904 38304
rect 85456 38056 85568 38136
rect 85456 38000 85484 38056
rect 85540 38000 85568 38056
rect 85456 36819 85568 38000
rect 85456 36763 85482 36819
rect 85538 36763 85568 36819
rect 85456 36736 85568 36763
rect 85624 37716 85736 37800
rect 85624 37660 85653 37716
rect 85709 37660 85736 37716
rect 85624 36820 85736 37660
rect 85624 36764 85655 36820
rect 85711 36764 85736 36820
rect 85624 36736 85736 36764
rect 91112 37381 91224 37464
rect 91112 37325 91140 37381
rect 91196 37325 91224 37381
rect 91112 36821 91224 37325
rect 91280 37408 92456 37464
rect 91280 37296 91366 37408
rect 91478 37296 92232 37408
rect 92344 37296 92456 37408
rect 91280 37240 92456 37296
rect 91112 36765 91140 36821
rect 91196 36765 91224 36821
rect 91112 36736 91224 36765
rect 87696 35481 87808 35486
rect 87696 35425 87716 35481
rect 87772 35425 87808 35481
rect 85176 35336 86288 35392
rect 85176 35280 86222 35336
rect 86278 35280 86288 35336
rect 85176 35224 86288 35280
rect 84748 34802 84860 34888
rect 84748 34746 84779 34802
rect 84835 34746 84860 34802
rect 84748 34664 84860 34746
rect 81368 34413 81397 34469
rect 81453 34413 81480 34469
rect 81368 34328 81480 34413
rect 79128 33179 79154 33235
rect 79210 33179 79240 33235
rect 79128 33152 79240 33179
rect 79296 34132 79408 34216
rect 79296 34076 79325 34132
rect 79381 34076 79408 34132
rect 79296 33231 79408 34076
rect 79296 33175 79331 33231
rect 79387 33175 79408 33231
rect 79296 33152 79408 33175
rect 84784 33797 84896 33880
rect 84784 33741 84812 33797
rect 84868 33741 84896 33797
rect 84784 33237 84896 33741
rect 84784 33181 84812 33237
rect 84868 33181 84896 33237
rect 84784 33152 84896 33181
rect 81368 31897 81480 31902
rect 81368 31841 81388 31897
rect 81444 31841 81480 31897
rect 78848 31752 79960 31808
rect 78848 31696 79894 31752
rect 79950 31696 79960 31752
rect 78848 31640 79960 31696
rect 78420 31218 78532 31304
rect 78420 31162 78451 31218
rect 78507 31162 78532 31218
rect 78420 31080 78532 31162
rect 75040 30829 75069 30885
rect 75125 30829 75152 30885
rect 75040 30744 75152 30829
rect 72800 29594 72824 29650
rect 72880 29594 72912 29650
rect 72800 29568 72912 29594
rect 72968 30548 73080 30632
rect 72968 30492 72997 30548
rect 73053 30492 73080 30548
rect 72968 29651 73080 30492
rect 72968 29595 72995 29651
rect 73051 29595 73080 29651
rect 72968 29568 73080 29595
rect 78456 30213 78568 30296
rect 78456 30157 78484 30213
rect 78540 30157 78568 30213
rect 78456 29653 78568 30157
rect 78456 29597 78484 29653
rect 78540 29597 78568 29653
rect 78456 29568 78568 29597
rect 75040 28313 75152 28318
rect 75040 28257 75060 28313
rect 75116 28257 75152 28313
rect 72520 28168 73632 28224
rect 72520 28112 73566 28168
rect 73622 28112 73632 28168
rect 72520 28056 73632 28112
rect 72092 27634 72204 27720
rect 72092 27578 72123 27634
rect 72179 27578 72204 27634
rect 72092 27496 72204 27578
rect 68712 27245 68741 27301
rect 68797 27245 68824 27301
rect 68712 27160 68824 27245
rect 66472 26010 66499 26066
rect 66555 26010 66584 26066
rect 66472 25984 66584 26010
rect 66640 26964 66752 27048
rect 66640 26908 66669 26964
rect 66725 26908 66752 26964
rect 66640 26071 66752 26908
rect 66640 26015 66670 26071
rect 66726 26015 66752 26071
rect 66640 25984 66752 26015
rect 72128 26629 72240 26712
rect 72128 26573 72156 26629
rect 72212 26573 72240 26629
rect 72128 26069 72240 26573
rect 72128 26013 72156 26069
rect 72212 26013 72240 26069
rect 72128 25984 72240 26013
rect 68712 24729 68824 24734
rect 68712 24673 68732 24729
rect 68788 24673 68824 24729
rect 66192 24584 67304 24640
rect 66192 24528 67238 24584
rect 67294 24528 67304 24584
rect 66192 24472 67304 24528
rect 65764 24050 65876 24136
rect 65764 23994 65795 24050
rect 65851 23994 65876 24050
rect 65764 23912 65876 23994
rect 62384 23661 62413 23717
rect 62469 23661 62496 23717
rect 62384 23576 62496 23661
rect 60144 22423 60164 22479
rect 60220 22423 60256 22479
rect 60144 22400 60256 22423
rect 60312 23380 60424 23464
rect 60312 23324 60341 23380
rect 60397 23324 60424 23380
rect 60312 22488 60424 23324
rect 60312 22432 60339 22488
rect 60395 22432 60424 22488
rect 60312 22400 60424 22432
rect 65800 23045 65912 23128
rect 65800 22989 65828 23045
rect 65884 22989 65912 23045
rect 65800 22485 65912 22989
rect 65800 22429 65828 22485
rect 65884 22429 65912 22485
rect 65800 22400 65912 22429
rect 62384 21145 62496 21150
rect 62384 21089 62404 21145
rect 62460 21089 62496 21145
rect 59864 21000 60976 21056
rect 59864 20944 60910 21000
rect 60966 20944 60976 21000
rect 59864 20888 60976 20944
rect 59436 20466 59548 20552
rect 59436 20410 59467 20466
rect 59523 20410 59548 20466
rect 59436 20328 59548 20410
rect 56056 20077 56085 20133
rect 56141 20077 56168 20133
rect 56056 19992 56168 20077
rect 53816 18847 53847 18903
rect 53903 18847 53928 18903
rect 53816 18816 53928 18847
rect 53984 19796 54096 19880
rect 53984 19740 54013 19796
rect 54069 19740 54096 19796
rect 53984 18899 54096 19740
rect 53984 18843 54010 18899
rect 54066 18843 54096 18899
rect 53984 18816 54096 18843
rect 59472 19461 59584 19544
rect 59472 19405 59500 19461
rect 59556 19405 59584 19461
rect 59472 18901 59584 19405
rect 59472 18845 59500 18901
rect 59556 18845 59584 18901
rect 59472 18816 59584 18845
rect 56056 17561 56168 17566
rect 56056 17505 56076 17561
rect 56132 17505 56168 17561
rect 53536 17416 54648 17472
rect 53536 17360 54582 17416
rect 54638 17360 54648 17416
rect 53536 17304 54648 17360
rect 53108 16882 53220 16968
rect 53108 16826 53139 16882
rect 53195 16826 53220 16882
rect 53108 16744 53220 16826
rect 49728 16493 49757 16549
rect 49813 16493 49840 16549
rect 49728 16408 49840 16493
rect 47488 15258 47514 15314
rect 47570 15258 47600 15314
rect 47488 15232 47600 15258
rect 47656 16212 47768 16296
rect 47656 16156 47685 16212
rect 47741 16156 47768 16212
rect 47656 15316 47768 16156
rect 47656 15260 47683 15316
rect 47739 15260 47768 15316
rect 47656 15232 47768 15260
rect 53144 15877 53256 15960
rect 53144 15821 53172 15877
rect 53228 15821 53256 15877
rect 53144 15317 53256 15821
rect 53144 15261 53172 15317
rect 53228 15261 53256 15317
rect 53144 15232 53256 15261
rect 49728 13977 49840 13982
rect 49728 13921 49748 13977
rect 49804 13921 49840 13977
rect 47208 13832 48320 13888
rect 47208 13776 48254 13832
rect 48310 13776 48320 13832
rect 47208 13720 48320 13776
rect 46780 13298 46892 13384
rect 46780 13242 46811 13298
rect 46867 13242 46892 13298
rect 46780 13160 46892 13242
rect 43400 12909 43429 12965
rect 43485 12909 43512 12965
rect 43400 12824 43512 12909
rect 44379 12992 44723 13048
rect 44379 12880 44497 12992
rect 44609 12880 44723 12992
rect 44379 12824 44723 12880
rect 47208 12656 47376 13720
rect 47959 12992 48303 13048
rect 47959 12880 48071 12992
rect 48183 12880 48303 12992
rect 47959 12824 48303 12880
rect 49250 12992 49594 13048
rect 49250 12880 49364 12992
rect 49476 12880 49594 12992
rect 49250 12824 49594 12880
rect 49728 12965 49840 13921
rect 53125 13384 53201 14056
rect 53536 13888 53704 17304
rect 53816 16552 53928 16632
rect 53816 16496 53844 16552
rect 53900 16496 53928 16552
rect 53816 15314 53928 16496
rect 56056 16549 56168 17505
rect 59453 16968 59529 17640
rect 59864 17472 60032 20888
rect 60144 20136 60256 20216
rect 60144 20080 60172 20136
rect 60228 20080 60256 20136
rect 60144 18898 60256 20080
rect 62384 20133 62496 21089
rect 65781 20552 65857 21224
rect 66192 21056 66360 24472
rect 66472 23720 66584 23800
rect 66472 23664 66500 23720
rect 66556 23664 66584 23720
rect 66472 22483 66584 23664
rect 68712 23717 68824 24673
rect 72109 24136 72185 24808
rect 72520 24640 72688 28056
rect 72800 27304 72912 27384
rect 72800 27248 72828 27304
rect 72884 27248 72912 27304
rect 72800 26068 72912 27248
rect 75040 27301 75152 28257
rect 78437 27720 78513 28392
rect 78848 28224 79016 31640
rect 79128 30888 79240 30968
rect 79128 30832 79156 30888
rect 79212 30832 79240 30888
rect 79128 29648 79240 30832
rect 81368 30885 81480 31841
rect 84765 31304 84841 31976
rect 85176 31808 85344 35224
rect 85456 34472 85568 34552
rect 85456 34416 85484 34472
rect 85540 34416 85568 34472
rect 85456 33233 85568 34416
rect 87696 34469 87808 35425
rect 91093 34888 91169 35560
rect 91076 34802 91188 34888
rect 91076 34746 91107 34802
rect 91163 34746 91188 34802
rect 91076 34664 91188 34746
rect 91280 34832 92904 34888
rect 91280 34720 91360 34832
rect 91472 34720 92680 34832
rect 92792 34720 92904 34832
rect 91280 34664 92904 34720
rect 87696 34413 87725 34469
rect 87781 34413 87808 34469
rect 87696 34328 87808 34413
rect 85456 33177 85479 33233
rect 85535 33177 85568 33233
rect 85456 33152 85568 33177
rect 85624 34132 85736 34216
rect 85624 34076 85653 34132
rect 85709 34076 85736 34132
rect 85624 33235 85736 34076
rect 85624 33179 85652 33235
rect 85708 33179 85736 33235
rect 85624 33152 85736 33179
rect 91112 33797 91224 33880
rect 91112 33741 91140 33797
rect 91196 33741 91224 33797
rect 91112 33237 91224 33741
rect 91280 33824 92456 33880
rect 91280 33712 91359 33824
rect 91471 33712 92232 33824
rect 92344 33712 92456 33824
rect 91280 33656 92456 33712
rect 91112 33181 91140 33237
rect 91196 33181 91224 33237
rect 91112 33152 91224 33181
rect 87696 31897 87808 31902
rect 87696 31841 87716 31897
rect 87772 31841 87808 31897
rect 85176 31752 86288 31808
rect 85176 31696 86222 31752
rect 86278 31696 86288 31752
rect 85176 31640 86288 31696
rect 84748 31218 84860 31304
rect 84748 31162 84779 31218
rect 84835 31162 84860 31218
rect 84748 31080 84860 31162
rect 81368 30829 81397 30885
rect 81453 30829 81480 30885
rect 81368 30744 81480 30829
rect 79128 29592 79149 29648
rect 79205 29592 79240 29648
rect 79128 29568 79240 29592
rect 79296 30548 79408 30632
rect 79296 30492 79325 30548
rect 79381 30492 79408 30548
rect 79296 29652 79408 30492
rect 79296 29596 79323 29652
rect 79379 29596 79408 29652
rect 79296 29568 79408 29596
rect 84784 30213 84896 30296
rect 84784 30157 84812 30213
rect 84868 30157 84896 30213
rect 84784 29653 84896 30157
rect 84784 29597 84812 29653
rect 84868 29597 84896 29653
rect 84784 29568 84896 29597
rect 81368 28313 81480 28318
rect 81368 28257 81388 28313
rect 81444 28257 81480 28313
rect 78848 28168 79960 28224
rect 78848 28112 79894 28168
rect 79950 28112 79960 28168
rect 78848 28056 79960 28112
rect 78420 27634 78532 27720
rect 78420 27578 78451 27634
rect 78507 27578 78532 27634
rect 78420 27496 78532 27578
rect 75040 27245 75069 27301
rect 75125 27245 75152 27301
rect 75040 27160 75152 27245
rect 72800 26012 72829 26068
rect 72885 26012 72912 26068
rect 72800 25984 72912 26012
rect 72968 26964 73080 27048
rect 72968 26908 72997 26964
rect 73053 26908 73080 26964
rect 72968 26067 73080 26908
rect 72968 26011 72998 26067
rect 73054 26011 73080 26067
rect 72968 25984 73080 26011
rect 78456 26629 78568 26712
rect 78456 26573 78484 26629
rect 78540 26573 78568 26629
rect 78456 26069 78568 26573
rect 78456 26013 78484 26069
rect 78540 26013 78568 26069
rect 78456 25984 78568 26013
rect 75040 24729 75152 24734
rect 75040 24673 75060 24729
rect 75116 24673 75152 24729
rect 72520 24584 73632 24640
rect 72520 24528 73566 24584
rect 73622 24528 73632 24584
rect 72520 24472 73632 24528
rect 72092 24050 72204 24136
rect 72092 23994 72123 24050
rect 72179 23994 72204 24050
rect 72092 23912 72204 23994
rect 68712 23661 68741 23717
rect 68797 23661 68824 23717
rect 68712 23576 68824 23661
rect 66472 22427 66498 22483
rect 66554 22427 66584 22483
rect 66472 22400 66584 22427
rect 66640 23380 66752 23464
rect 66640 23324 66669 23380
rect 66725 23324 66752 23380
rect 66640 22488 66752 23324
rect 66640 22432 66666 22488
rect 66722 22432 66752 22488
rect 66640 22400 66752 22432
rect 72128 23045 72240 23128
rect 72128 22989 72156 23045
rect 72212 22989 72240 23045
rect 72128 22485 72240 22989
rect 72128 22429 72156 22485
rect 72212 22429 72240 22485
rect 72128 22400 72240 22429
rect 68712 21145 68824 21150
rect 68712 21089 68732 21145
rect 68788 21089 68824 21145
rect 66192 21000 67304 21056
rect 66192 20944 67238 21000
rect 67294 20944 67304 21000
rect 66192 20888 67304 20944
rect 65764 20466 65876 20552
rect 65764 20410 65795 20466
rect 65851 20410 65876 20466
rect 65764 20328 65876 20410
rect 62384 20077 62413 20133
rect 62469 20077 62496 20133
rect 62384 19992 62496 20077
rect 60144 18842 60174 18898
rect 60230 18842 60256 18898
rect 60144 18816 60256 18842
rect 60312 19796 60424 19880
rect 60312 19740 60341 19796
rect 60397 19740 60424 19796
rect 60312 18898 60424 19740
rect 60312 18842 60339 18898
rect 60395 18842 60424 18898
rect 60312 18816 60424 18842
rect 65800 19461 65912 19544
rect 65800 19405 65828 19461
rect 65884 19405 65912 19461
rect 65800 18901 65912 19405
rect 65800 18845 65828 18901
rect 65884 18845 65912 18901
rect 65800 18816 65912 18845
rect 62384 17561 62496 17566
rect 62384 17505 62404 17561
rect 62460 17505 62496 17561
rect 59864 17416 60976 17472
rect 59864 17360 60910 17416
rect 60966 17360 60976 17416
rect 59864 17304 60976 17360
rect 59436 16882 59548 16968
rect 59436 16826 59467 16882
rect 59523 16826 59548 16882
rect 59436 16744 59548 16826
rect 56056 16493 56085 16549
rect 56141 16493 56168 16549
rect 56056 16408 56168 16493
rect 53816 15258 53842 15314
rect 53898 15258 53928 15314
rect 53816 15232 53928 15258
rect 53984 16212 54096 16296
rect 53984 16156 54013 16212
rect 54069 16156 54096 16212
rect 53984 15316 54096 16156
rect 53984 15260 54013 15316
rect 54069 15260 54096 15316
rect 53984 15232 54096 15260
rect 59472 15877 59584 15960
rect 59472 15821 59500 15877
rect 59556 15821 59584 15877
rect 59472 15317 59584 15821
rect 59472 15261 59500 15317
rect 59556 15261 59584 15317
rect 59472 15232 59584 15261
rect 56056 13977 56168 13982
rect 56056 13921 56076 13977
rect 56132 13921 56168 13977
rect 53536 13832 54648 13888
rect 53536 13776 54582 13832
rect 54638 13776 54648 13832
rect 53536 13720 54648 13776
rect 53108 13298 53220 13384
rect 53108 13242 53139 13298
rect 53195 13242 53220 13298
rect 53108 13160 53220 13242
rect 49728 12909 49757 12965
rect 49813 12909 49840 12965
rect 49728 12824 49840 12909
rect 50707 12992 51051 13048
rect 50707 12880 50820 12992
rect 50932 12880 51051 12992
rect 50707 12824 51051 12880
rect 53536 12656 53704 13720
rect 54286 12992 54630 13048
rect 54286 12880 54399 12992
rect 54511 12880 54630 12992
rect 54286 12824 54630 12880
rect 55578 12992 55922 13048
rect 55578 12880 55689 12992
rect 55801 12880 55922 12992
rect 55578 12824 55922 12880
rect 56056 12965 56168 13921
rect 59453 13384 59529 14056
rect 59864 13888 60032 17304
rect 60144 16552 60256 16632
rect 60144 16496 60172 16552
rect 60228 16496 60256 16552
rect 60144 15309 60256 16496
rect 62384 16549 62496 17505
rect 65781 16968 65857 17640
rect 66192 17472 66360 20888
rect 66472 20136 66584 20216
rect 66472 20080 66500 20136
rect 66556 20080 66584 20136
rect 66472 18900 66584 20080
rect 68712 20133 68824 21089
rect 72109 20552 72185 21224
rect 72520 21056 72688 24472
rect 72800 23720 72912 23800
rect 72800 23664 72828 23720
rect 72884 23664 72912 23720
rect 72800 22487 72912 23664
rect 75040 23717 75152 24673
rect 78437 24136 78513 24808
rect 78848 24640 79016 28056
rect 79128 27304 79240 27384
rect 79128 27248 79156 27304
rect 79212 27248 79240 27304
rect 79128 26071 79240 27248
rect 81368 27301 81480 28257
rect 84765 27720 84841 28392
rect 85176 28224 85344 31640
rect 85456 30888 85568 30968
rect 85456 30832 85484 30888
rect 85540 30832 85568 30888
rect 85456 29652 85568 30832
rect 87696 30885 87808 31841
rect 91093 31304 91169 31976
rect 91076 31218 91188 31304
rect 91076 31162 91107 31218
rect 91163 31162 91188 31218
rect 91076 31080 91188 31162
rect 91280 31248 92904 31304
rect 91280 31136 91362 31248
rect 91474 31136 92680 31248
rect 92792 31136 92904 31248
rect 91280 31080 92904 31136
rect 87696 30829 87725 30885
rect 87781 30829 87808 30885
rect 87696 30744 87808 30829
rect 85456 29596 85483 29652
rect 85539 29596 85568 29652
rect 85456 29568 85568 29596
rect 85624 30548 85736 30632
rect 85624 30492 85653 30548
rect 85709 30492 85736 30548
rect 85624 29650 85736 30492
rect 85624 29594 85659 29650
rect 85715 29594 85736 29650
rect 85624 29568 85736 29594
rect 91112 30213 91224 30296
rect 91112 30157 91140 30213
rect 91196 30157 91224 30213
rect 91112 29653 91224 30157
rect 91280 30240 92456 30296
rect 91280 30128 91365 30240
rect 91477 30128 92232 30240
rect 92344 30128 92456 30240
rect 91280 30072 92456 30128
rect 91112 29597 91140 29653
rect 91196 29597 91224 29653
rect 91112 29568 91224 29597
rect 87696 28313 87808 28318
rect 87696 28257 87716 28313
rect 87772 28257 87808 28313
rect 85176 28168 86288 28224
rect 85176 28112 86222 28168
rect 86278 28112 86288 28168
rect 85176 28056 86288 28112
rect 84748 27634 84860 27720
rect 84748 27578 84779 27634
rect 84835 27578 84860 27634
rect 84748 27496 84860 27578
rect 81368 27245 81397 27301
rect 81453 27245 81480 27301
rect 81368 27160 81480 27245
rect 79128 26015 79156 26071
rect 79212 26015 79240 26071
rect 79128 25984 79240 26015
rect 79296 26964 79408 27048
rect 79296 26908 79325 26964
rect 79381 26908 79408 26964
rect 79296 26066 79408 26908
rect 79296 26010 79325 26066
rect 79381 26010 79408 26066
rect 79296 25984 79408 26010
rect 84784 26629 84896 26712
rect 84784 26573 84812 26629
rect 84868 26573 84896 26629
rect 84784 26069 84896 26573
rect 84784 26013 84812 26069
rect 84868 26013 84896 26069
rect 84784 25984 84896 26013
rect 81368 24729 81480 24734
rect 81368 24673 81388 24729
rect 81444 24673 81480 24729
rect 78848 24584 79960 24640
rect 78848 24528 79894 24584
rect 79950 24528 79960 24584
rect 78848 24472 79960 24528
rect 78420 24050 78532 24136
rect 78420 23994 78451 24050
rect 78507 23994 78532 24050
rect 78420 23912 78532 23994
rect 75040 23661 75069 23717
rect 75125 23661 75152 23717
rect 75040 23576 75152 23661
rect 72800 22431 72832 22487
rect 72888 22431 72912 22487
rect 72800 22400 72912 22431
rect 72968 23380 73080 23464
rect 72968 23324 72997 23380
rect 73053 23324 73080 23380
rect 72968 22483 73080 23324
rect 72968 22427 72989 22483
rect 73045 22427 73080 22483
rect 72968 22400 73080 22427
rect 78456 23045 78568 23128
rect 78456 22989 78484 23045
rect 78540 22989 78568 23045
rect 78456 22485 78568 22989
rect 78456 22429 78484 22485
rect 78540 22429 78568 22485
rect 78456 22400 78568 22429
rect 75040 21145 75152 21150
rect 75040 21089 75060 21145
rect 75116 21089 75152 21145
rect 72520 21000 73632 21056
rect 72520 20944 73566 21000
rect 73622 20944 73632 21000
rect 72520 20888 73632 20944
rect 72092 20466 72204 20552
rect 72092 20410 72123 20466
rect 72179 20410 72204 20466
rect 72092 20328 72204 20410
rect 68712 20077 68741 20133
rect 68797 20077 68824 20133
rect 68712 19992 68824 20077
rect 66472 18844 66500 18900
rect 66556 18844 66584 18900
rect 66472 18816 66584 18844
rect 66640 19796 66752 19880
rect 66640 19740 66669 19796
rect 66725 19740 66752 19796
rect 66640 18899 66752 19740
rect 66640 18843 66667 18899
rect 66723 18843 66752 18899
rect 66640 18816 66752 18843
rect 72128 19461 72240 19544
rect 72128 19405 72156 19461
rect 72212 19405 72240 19461
rect 72128 18901 72240 19405
rect 72128 18845 72156 18901
rect 72212 18845 72240 18901
rect 72128 18816 72240 18845
rect 68712 17561 68824 17566
rect 68712 17505 68732 17561
rect 68788 17505 68824 17561
rect 66192 17416 67304 17472
rect 66192 17360 67238 17416
rect 67294 17360 67304 17416
rect 66192 17304 67304 17360
rect 65764 16882 65876 16968
rect 65764 16826 65795 16882
rect 65851 16826 65876 16882
rect 65764 16744 65876 16826
rect 62384 16493 62413 16549
rect 62469 16493 62496 16549
rect 62384 16408 62496 16493
rect 60144 15253 60166 15309
rect 60222 15253 60256 15309
rect 60144 15232 60256 15253
rect 60312 16212 60424 16296
rect 60312 16156 60341 16212
rect 60397 16156 60424 16212
rect 60312 15314 60424 16156
rect 60312 15258 60343 15314
rect 60399 15258 60424 15314
rect 60312 15232 60424 15258
rect 65800 15877 65912 15960
rect 65800 15821 65828 15877
rect 65884 15821 65912 15877
rect 65800 15317 65912 15821
rect 65800 15261 65828 15317
rect 65884 15261 65912 15317
rect 65800 15232 65912 15261
rect 62384 13977 62496 13982
rect 62384 13921 62404 13977
rect 62460 13921 62496 13977
rect 59864 13832 60976 13888
rect 59864 13776 60910 13832
rect 60966 13776 60976 13832
rect 59864 13720 60976 13776
rect 59436 13298 59548 13384
rect 59436 13242 59467 13298
rect 59523 13242 59548 13298
rect 59436 13160 59548 13242
rect 56056 12909 56085 12965
rect 56141 12909 56168 12965
rect 56056 12824 56168 12909
rect 57035 12992 57379 13048
rect 57035 12880 57144 12992
rect 57256 12880 57379 12992
rect 57035 12824 57379 12880
rect 59864 12656 60032 13720
rect 60614 12824 60958 13048
rect 61906 12824 62250 13048
rect 62384 12965 62496 13921
rect 65781 13384 65857 14056
rect 66192 13888 66360 17304
rect 66472 16552 66584 16632
rect 66472 16496 66500 16552
rect 66556 16496 66584 16552
rect 66472 15315 66584 16496
rect 68712 16549 68824 17505
rect 72109 16968 72185 17640
rect 72520 17472 72688 20888
rect 72800 20136 72912 20216
rect 72800 20080 72828 20136
rect 72884 20080 72912 20136
rect 72800 18899 72912 20080
rect 75040 20133 75152 21089
rect 78437 20552 78513 21224
rect 78848 21056 79016 24472
rect 79128 23720 79240 23800
rect 79128 23664 79156 23720
rect 79212 23664 79240 23720
rect 79128 22480 79240 23664
rect 81368 23717 81480 24673
rect 84765 24136 84841 24808
rect 85176 24640 85344 28056
rect 85456 27304 85568 27384
rect 85456 27248 85484 27304
rect 85540 27248 85568 27304
rect 85456 26071 85568 27248
rect 87696 27301 87808 28257
rect 91093 27720 91169 28392
rect 91076 27634 91188 27720
rect 91076 27578 91107 27634
rect 91163 27578 91188 27634
rect 91076 27496 91188 27578
rect 91280 27664 92904 27720
rect 91280 27552 91364 27664
rect 91476 27552 92680 27664
rect 92792 27552 92904 27664
rect 91280 27496 92904 27552
rect 87696 27245 87725 27301
rect 87781 27245 87808 27301
rect 87696 27160 87808 27245
rect 85456 26015 85486 26071
rect 85542 26015 85568 26071
rect 85456 25984 85568 26015
rect 85624 26964 85736 27048
rect 85624 26908 85653 26964
rect 85709 26908 85736 26964
rect 85624 26068 85736 26908
rect 85624 26012 85655 26068
rect 85711 26012 85736 26068
rect 85624 25984 85736 26012
rect 91112 26629 91224 26712
rect 91112 26573 91140 26629
rect 91196 26573 91224 26629
rect 91112 26069 91224 26573
rect 91280 26656 92456 26712
rect 91280 26544 91364 26656
rect 91476 26544 92232 26656
rect 92344 26544 92456 26656
rect 91280 26488 92456 26544
rect 91112 26013 91140 26069
rect 91196 26013 91224 26069
rect 91112 25984 91224 26013
rect 87696 24729 87808 24734
rect 87696 24673 87716 24729
rect 87772 24673 87808 24729
rect 85176 24584 86288 24640
rect 85176 24528 86222 24584
rect 86278 24528 86288 24584
rect 85176 24472 86288 24528
rect 84748 24050 84860 24136
rect 84748 23994 84779 24050
rect 84835 23994 84860 24050
rect 84748 23912 84860 23994
rect 81368 23661 81397 23717
rect 81453 23661 81480 23717
rect 81368 23576 81480 23661
rect 79128 22424 79152 22480
rect 79208 22424 79240 22480
rect 79128 22400 79240 22424
rect 79296 23380 79408 23464
rect 79296 23324 79325 23380
rect 79381 23324 79408 23380
rect 79296 22483 79408 23324
rect 79296 22427 79323 22483
rect 79379 22427 79408 22483
rect 79296 22400 79408 22427
rect 84784 23045 84896 23128
rect 84784 22989 84812 23045
rect 84868 22989 84896 23045
rect 84784 22485 84896 22989
rect 84784 22429 84812 22485
rect 84868 22429 84896 22485
rect 84784 22400 84896 22429
rect 81368 21145 81480 21150
rect 81368 21089 81388 21145
rect 81444 21089 81480 21145
rect 78848 21000 79960 21056
rect 78848 20944 79894 21000
rect 79950 20944 79960 21000
rect 78848 20888 79960 20944
rect 78420 20466 78532 20552
rect 78420 20410 78451 20466
rect 78507 20410 78532 20466
rect 78420 20328 78532 20410
rect 75040 20077 75069 20133
rect 75125 20077 75152 20133
rect 75040 19992 75152 20077
rect 72800 18843 72830 18899
rect 72886 18843 72912 18899
rect 72800 18816 72912 18843
rect 72968 19796 73080 19880
rect 72968 19740 72997 19796
rect 73053 19740 73080 19796
rect 72968 18899 73080 19740
rect 72968 18843 72999 18899
rect 73055 18843 73080 18899
rect 72968 18816 73080 18843
rect 78456 19461 78568 19544
rect 78456 19405 78484 19461
rect 78540 19405 78568 19461
rect 78456 18901 78568 19405
rect 78456 18845 78484 18901
rect 78540 18845 78568 18901
rect 78456 18816 78568 18845
rect 75040 17561 75152 17566
rect 75040 17505 75060 17561
rect 75116 17505 75152 17561
rect 72520 17416 73632 17472
rect 72520 17360 73566 17416
rect 73622 17360 73632 17416
rect 72520 17304 73632 17360
rect 72092 16882 72204 16968
rect 72092 16826 72123 16882
rect 72179 16826 72204 16882
rect 72092 16744 72204 16826
rect 68712 16493 68741 16549
rect 68797 16493 68824 16549
rect 68712 16408 68824 16493
rect 66472 15259 66498 15315
rect 66554 15259 66584 15315
rect 66472 15232 66584 15259
rect 66640 16212 66752 16296
rect 66640 16156 66669 16212
rect 66725 16156 66752 16212
rect 66640 15316 66752 16156
rect 66640 15260 66665 15316
rect 66721 15260 66752 15316
rect 66640 15232 66752 15260
rect 72128 15877 72240 15960
rect 72128 15821 72156 15877
rect 72212 15821 72240 15877
rect 72128 15317 72240 15821
rect 72128 15261 72156 15317
rect 72212 15261 72240 15317
rect 72128 15232 72240 15261
rect 68712 13977 68824 13982
rect 68712 13921 68732 13977
rect 68788 13921 68824 13977
rect 66192 13832 67304 13888
rect 66192 13776 67238 13832
rect 67294 13776 67304 13832
rect 66192 13720 67304 13776
rect 65764 13298 65876 13384
rect 65764 13242 65795 13298
rect 65851 13242 65876 13298
rect 65764 13160 65876 13242
rect 62384 12909 62413 12965
rect 62469 12909 62496 12965
rect 62384 12824 62496 12909
rect 63363 12824 63707 13048
rect 66192 12656 66360 13720
rect 66942 12824 67286 13048
rect 68234 12824 68578 13048
rect 68712 12965 68824 13921
rect 72109 13384 72185 14056
rect 72520 13888 72688 17304
rect 72800 16552 72912 16632
rect 72800 16496 72828 16552
rect 72884 16496 72912 16552
rect 72800 15318 72912 16496
rect 75040 16549 75152 17505
rect 78437 16968 78513 17640
rect 78848 17472 79016 20888
rect 79128 20136 79240 20216
rect 79128 20080 79156 20136
rect 79212 20080 79240 20136
rect 79128 18901 79240 20080
rect 81368 20133 81480 21089
rect 84765 20552 84841 21224
rect 85176 21056 85344 24472
rect 85456 23720 85568 23800
rect 85456 23664 85484 23720
rect 85540 23664 85568 23720
rect 85456 22480 85568 23664
rect 87696 23717 87808 24673
rect 91093 24136 91169 24808
rect 91076 24050 91188 24136
rect 91076 23994 91107 24050
rect 91163 23994 91188 24050
rect 91076 23912 91188 23994
rect 91280 24080 92904 24136
rect 91280 23968 91365 24080
rect 91477 23968 92680 24080
rect 92792 23968 92904 24080
rect 91280 23912 92904 23968
rect 87696 23661 87725 23717
rect 87781 23661 87808 23717
rect 87696 23576 87808 23661
rect 85456 22424 85481 22480
rect 85537 22424 85568 22480
rect 85456 22400 85568 22424
rect 85624 23380 85736 23464
rect 85624 23324 85653 23380
rect 85709 23324 85736 23380
rect 85624 22482 85736 23324
rect 85624 22426 85655 22482
rect 85711 22426 85736 22482
rect 85624 22400 85736 22426
rect 91112 23045 91224 23128
rect 91112 22989 91140 23045
rect 91196 22989 91224 23045
rect 91112 22485 91224 22989
rect 91280 23072 92456 23128
rect 91280 22960 91363 23072
rect 91475 22960 92232 23072
rect 92344 22960 92456 23072
rect 91280 22904 92456 22960
rect 91112 22429 91140 22485
rect 91196 22429 91224 22485
rect 91112 22400 91224 22429
rect 87696 21145 87808 21150
rect 87696 21089 87716 21145
rect 87772 21089 87808 21145
rect 85176 21000 86288 21056
rect 85176 20944 86222 21000
rect 86278 20944 86288 21000
rect 85176 20888 86288 20944
rect 84748 20466 84860 20552
rect 84748 20410 84779 20466
rect 84835 20410 84860 20466
rect 84748 20328 84860 20410
rect 81368 20077 81397 20133
rect 81453 20077 81480 20133
rect 81368 19992 81480 20077
rect 79128 18845 79159 18901
rect 79215 18845 79240 18901
rect 79128 18816 79240 18845
rect 79296 19796 79408 19880
rect 79296 19740 79325 19796
rect 79381 19740 79408 19796
rect 79296 18900 79408 19740
rect 79296 18844 79327 18900
rect 79383 18844 79408 18900
rect 79296 18816 79408 18844
rect 84784 19461 84896 19544
rect 84784 19405 84812 19461
rect 84868 19405 84896 19461
rect 84784 18901 84896 19405
rect 84784 18845 84812 18901
rect 84868 18845 84896 18901
rect 84784 18816 84896 18845
rect 81368 17561 81480 17566
rect 81368 17505 81388 17561
rect 81444 17505 81480 17561
rect 78848 17416 79960 17472
rect 78848 17360 79894 17416
rect 79950 17360 79960 17416
rect 78848 17304 79960 17360
rect 78420 16882 78532 16968
rect 78420 16826 78451 16882
rect 78507 16826 78532 16882
rect 78420 16744 78532 16826
rect 75040 16493 75069 16549
rect 75125 16493 75152 16549
rect 75040 16408 75152 16493
rect 72800 15262 72829 15318
rect 72885 15262 72912 15318
rect 72800 15232 72912 15262
rect 72968 16212 73080 16296
rect 72968 16156 72997 16212
rect 73053 16156 73080 16212
rect 72968 15316 73080 16156
rect 72968 15260 72994 15316
rect 73050 15260 73080 15316
rect 72968 15232 73080 15260
rect 78456 15877 78568 15960
rect 78456 15821 78484 15877
rect 78540 15821 78568 15877
rect 78456 15317 78568 15821
rect 78456 15261 78484 15317
rect 78540 15261 78568 15317
rect 78456 15232 78568 15261
rect 75040 13977 75152 13982
rect 75040 13921 75060 13977
rect 75116 13921 75152 13977
rect 72520 13832 73632 13888
rect 72520 13776 73566 13832
rect 73622 13776 73632 13832
rect 72520 13720 73632 13776
rect 72092 13298 72204 13384
rect 72092 13242 72123 13298
rect 72179 13242 72204 13298
rect 72092 13160 72204 13242
rect 68712 12909 68741 12965
rect 68797 12909 68824 12965
rect 68712 12824 68824 12909
rect 69691 12824 70035 13048
rect 72520 12656 72688 13720
rect 73270 12824 73614 13048
rect 74562 12824 74906 13048
rect 75040 12965 75152 13921
rect 78437 13384 78513 14056
rect 78848 13888 79016 17304
rect 79128 16552 79240 16632
rect 79128 16496 79156 16552
rect 79212 16496 79240 16552
rect 79128 15314 79240 16496
rect 81368 16549 81480 17505
rect 84765 16968 84841 17640
rect 85176 17472 85344 20888
rect 85456 20136 85568 20216
rect 85456 20080 85484 20136
rect 85540 20080 85568 20136
rect 85456 18904 85568 20080
rect 87696 20133 87808 21089
rect 91093 20552 91169 21224
rect 91076 20466 91188 20552
rect 91076 20410 91107 20466
rect 91163 20410 91188 20466
rect 91076 20328 91188 20410
rect 91280 20496 92904 20552
rect 91280 20384 91363 20496
rect 91475 20384 92680 20496
rect 92792 20384 92904 20496
rect 91280 20328 92904 20384
rect 87696 20077 87725 20133
rect 87781 20077 87808 20133
rect 87696 19992 87808 20077
rect 85456 18848 85487 18904
rect 85543 18848 85568 18904
rect 85456 18816 85568 18848
rect 85624 19796 85736 19880
rect 85624 19740 85653 19796
rect 85709 19740 85736 19796
rect 85624 18899 85736 19740
rect 85624 18843 85651 18899
rect 85707 18843 85736 18899
rect 85624 18816 85736 18843
rect 91112 19461 91224 19544
rect 91112 19405 91140 19461
rect 91196 19405 91224 19461
rect 91112 18901 91224 19405
rect 91280 19488 92456 19544
rect 91280 19376 91365 19488
rect 91477 19376 92232 19488
rect 92344 19376 92456 19488
rect 91280 19320 92456 19376
rect 91112 18845 91140 18901
rect 91196 18845 91224 18901
rect 91112 18816 91224 18845
rect 87696 17561 87808 17566
rect 87696 17505 87716 17561
rect 87772 17505 87808 17561
rect 85176 17416 86288 17472
rect 85176 17360 86222 17416
rect 86278 17360 86288 17416
rect 85176 17304 86288 17360
rect 84748 16882 84860 16968
rect 84748 16826 84779 16882
rect 84835 16826 84860 16882
rect 84748 16744 84860 16826
rect 81368 16493 81397 16549
rect 81453 16493 81480 16549
rect 81368 16408 81480 16493
rect 79128 15258 79153 15314
rect 79209 15258 79240 15314
rect 79128 15232 79240 15258
rect 79296 16212 79408 16296
rect 79296 16156 79325 16212
rect 79381 16156 79408 16212
rect 79296 15313 79408 16156
rect 79296 15257 79325 15313
rect 79381 15257 79408 15313
rect 79296 15232 79408 15257
rect 84784 15877 84896 15960
rect 84784 15821 84812 15877
rect 84868 15821 84896 15877
rect 84784 15317 84896 15821
rect 84784 15261 84812 15317
rect 84868 15261 84896 15317
rect 84784 15232 84896 15261
rect 81368 13977 81480 13982
rect 81368 13921 81388 13977
rect 81444 13921 81480 13977
rect 78848 13832 79960 13888
rect 78848 13776 79894 13832
rect 79950 13776 79960 13832
rect 78848 13720 79960 13776
rect 78420 13298 78532 13384
rect 78420 13242 78451 13298
rect 78507 13242 78532 13298
rect 78420 13160 78532 13242
rect 75040 12909 75069 12965
rect 75125 12909 75152 12965
rect 75040 12824 75152 12909
rect 76019 12824 76363 13048
rect 78848 12656 79016 13720
rect 79598 12824 79942 13048
rect 80890 12824 81234 13048
rect 81368 12965 81480 13921
rect 84765 13384 84841 14056
rect 85176 13888 85344 17304
rect 85456 16552 85568 16632
rect 85456 16496 85484 16552
rect 85540 16496 85568 16552
rect 85456 15310 85568 16496
rect 87696 16549 87808 17505
rect 91093 16968 91169 17640
rect 91076 16882 91188 16968
rect 91076 16826 91107 16882
rect 91163 16826 91188 16882
rect 91076 16744 91188 16826
rect 91280 16912 92904 16968
rect 91280 16800 91362 16912
rect 91474 16800 92680 16912
rect 92792 16800 92904 16912
rect 91280 16744 92904 16800
rect 87696 16493 87725 16549
rect 87781 16493 87808 16549
rect 87696 16408 87808 16493
rect 85456 15254 85479 15310
rect 85535 15254 85568 15310
rect 85456 15232 85568 15254
rect 85624 16212 85736 16296
rect 85624 16156 85653 16212
rect 85709 16156 85736 16212
rect 85624 15314 85736 16156
rect 85624 15258 85649 15314
rect 85705 15258 85736 15314
rect 85624 15232 85736 15258
rect 91112 15877 91224 15960
rect 91112 15821 91140 15877
rect 91196 15821 91224 15877
rect 91112 15317 91224 15821
rect 91280 15904 92456 15960
rect 91280 15792 91356 15904
rect 91468 15792 92232 15904
rect 92344 15792 92456 15904
rect 91280 15736 92456 15792
rect 91112 15261 91140 15317
rect 91196 15261 91224 15317
rect 91112 15232 91224 15261
rect 87696 13977 87808 13982
rect 87696 13921 87716 13977
rect 87772 13921 87808 13977
rect 85176 13832 86288 13888
rect 85176 13776 86222 13832
rect 86278 13776 86288 13832
rect 85176 13720 86288 13776
rect 84748 13298 84860 13384
rect 84748 13242 84779 13298
rect 84835 13242 84860 13298
rect 84748 13160 84860 13242
rect 81368 12909 81397 12965
rect 81453 12909 81480 12965
rect 81368 12824 81480 12909
rect 82347 12824 82691 13048
rect 85176 12656 85344 13720
rect 85926 12824 86270 13048
rect 87218 12824 87562 13048
rect 87696 12965 87808 13921
rect 91093 13384 91169 14056
rect 91076 13298 91188 13384
rect 91076 13242 91107 13298
rect 91163 13242 91188 13298
rect 91076 13160 91188 13242
rect 91280 13328 92904 13384
rect 91280 13216 91366 13328
rect 91478 13216 92680 13328
rect 92792 13216 92904 13328
rect 91280 13160 92904 13216
rect 87696 12909 87725 12965
rect 87781 12909 87808 12965
rect 87696 12824 87808 12909
rect 88675 12824 89019 13048
<< via2 >>
rect 42392 41552 42504 41664
rect 43756 41552 43868 41664
rect 45212 41552 45324 41664
rect 48720 41552 48832 41664
rect 50088 41552 50200 41664
rect 51550 41552 51662 41664
rect 55048 41552 55160 41664
rect 56416 41552 56528 41664
rect 57873 41552 57985 41664
rect 61376 41552 61488 41664
rect 62746 41552 62858 41664
rect 64204 41552 64316 41664
rect 67704 41552 67816 41664
rect 69077 41552 69189 41664
rect 70528 41552 70640 41664
rect 74032 41552 74144 41664
rect 75403 41552 75515 41664
rect 76860 41552 76972 41664
rect 80360 41552 80472 41664
rect 81734 41552 81846 41664
rect 83186 41552 83298 41664
rect 41746 12880 41858 12992
rect 43036 12880 43148 12992
rect 44497 12880 44609 12992
rect 48071 12880 48183 12992
rect 49364 12880 49476 12992
rect 50820 12880 50932 12992
rect 54399 12880 54511 12992
rect 55689 12880 55801 12992
rect 57144 12880 57256 12992
<< metal3 >>
rect 42279 41664 42623 41719
rect 42279 41552 42392 41664
rect 42504 41552 42623 41664
rect 42279 41495 42623 41552
rect 43649 41664 43993 41720
rect 43649 41552 43756 41664
rect 43868 41552 43993 41664
rect 43649 41496 43993 41552
rect 45104 41664 45448 41720
rect 45104 41552 45212 41664
rect 45324 41552 45448 41664
rect 45104 41496 45448 41552
rect 48607 41664 48951 41720
rect 48607 41552 48720 41664
rect 48832 41552 48951 41664
rect 48607 41496 48951 41552
rect 49977 41664 50321 41720
rect 49977 41552 50088 41664
rect 50200 41552 50321 41664
rect 49977 41496 50321 41552
rect 51432 41664 51776 41720
rect 51432 41552 51550 41664
rect 51662 41552 51776 41664
rect 51432 41496 51776 41552
rect 54935 41664 55279 41720
rect 54935 41552 55048 41664
rect 55160 41552 55279 41664
rect 54935 41496 55279 41552
rect 56305 41664 56649 41720
rect 56305 41552 56416 41664
rect 56528 41552 56649 41664
rect 56305 41496 56649 41552
rect 57760 41664 58104 41720
rect 57760 41552 57873 41664
rect 57985 41552 58104 41664
rect 57760 41496 58104 41552
rect 61263 41664 61607 41720
rect 61263 41552 61376 41664
rect 61488 41552 61607 41664
rect 61263 41496 61607 41552
rect 62633 41664 62977 41720
rect 62633 41552 62746 41664
rect 62858 41552 62977 41664
rect 62633 41496 62977 41552
rect 64088 41664 64432 41720
rect 64088 41552 64204 41664
rect 64316 41552 64432 41664
rect 64088 41496 64432 41552
rect 67591 41664 67935 41720
rect 67591 41552 67704 41664
rect 67816 41552 67935 41664
rect 67591 41496 67935 41552
rect 68961 41664 69305 41720
rect 68961 41552 69077 41664
rect 69189 41552 69305 41664
rect 68961 41496 69305 41552
rect 70416 41664 70760 41720
rect 70416 41552 70528 41664
rect 70640 41552 70760 41664
rect 70416 41496 70760 41552
rect 73919 41664 74263 41720
rect 73919 41552 74032 41664
rect 74144 41552 74263 41664
rect 73919 41496 74263 41552
rect 75289 41664 75633 41720
rect 75289 41552 75403 41664
rect 75515 41552 75633 41664
rect 75289 41496 75633 41552
rect 76744 41664 77088 41720
rect 76744 41552 76860 41664
rect 76972 41552 77088 41664
rect 76744 41496 77088 41552
rect 80247 41664 80591 41720
rect 80247 41552 80360 41664
rect 80472 41552 80591 41664
rect 80247 41496 80591 41552
rect 81617 41664 81961 41720
rect 81617 41552 81734 41664
rect 81846 41552 81961 41664
rect 81617 41496 81961 41552
rect 83072 41664 83416 41720
rect 83072 41552 83186 41664
rect 83298 41552 83416 41664
rect 83072 41496 83416 41552
rect 41630 12992 41974 13048
rect 41630 12880 41746 12992
rect 41858 12880 41974 12992
rect 41630 12824 41974 12880
rect 42922 12992 43266 13048
rect 42922 12880 43036 12992
rect 43148 12880 43266 12992
rect 42922 12824 43266 12880
rect 44379 12992 44723 13048
rect 44379 12880 44497 12992
rect 44609 12880 44723 12992
rect 44379 12824 44723 12880
rect 47959 12992 48303 13048
rect 47959 12880 48071 12992
rect 48183 12880 48303 12992
rect 47959 12824 48303 12880
rect 49250 12992 49594 13048
rect 49250 12880 49364 12992
rect 49476 12880 49594 12992
rect 49250 12824 49594 12880
rect 50707 12992 51051 13048
rect 50707 12880 50820 12992
rect 50932 12880 51051 12992
rect 50707 12824 51051 12880
rect 54286 12992 54630 13048
rect 54286 12880 54399 12992
rect 54511 12880 54630 12992
rect 54286 12824 54630 12880
rect 55578 12992 55922 13048
rect 55578 12880 55689 12992
rect 55801 12880 55922 12992
rect 55578 12824 55922 12880
rect 57035 12992 57379 13048
rect 57035 12880 57144 12992
rect 57256 12880 57379 12992
rect 57035 12824 57379 12880
rect 60614 12824 60958 13048
rect 61906 12824 62250 13048
rect 63363 12824 63707 13048
rect 66942 12824 67286 13048
rect 68234 12824 68578 13048
rect 69691 12824 70035 13048
rect 73270 12824 73614 13048
rect 74562 12824 74906 13048
rect 76019 12824 76363 13048
rect 79598 12824 79942 13048
rect 80890 12824 81234 13048
rect 82347 12824 82691 13048
rect 85926 12824 86270 13048
rect 87218 12824 87562 13048
rect 88675 12824 89019 13048
<< metal4 >>
rect 66496 29592 66552 29648
rect 79149 29592 79205 29648
rect 85483 29596 85539 29652
use unit_cell_aray  unit_cell_aray_0
timestamp 1758523347
transform 1 0 85786 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_1
timestamp 1758523347
transform 1 0 79458 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_2
timestamp 1758523347
transform 1 0 73130 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_3
timestamp 1758523347
transform 1 0 66802 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_4
timestamp 1758523347
transform 1 0 54146 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_5
timestamp 1758523347
transform 1 0 60474 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_6
timestamp 1758523347
transform 1 0 47818 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_7
timestamp 1758523347
transform 1 0 41490 0 1 17321
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_8
timestamp 1758523347
transform 1 0 41490 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_9
timestamp 1758523347
transform 1 0 47818 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_10
timestamp 1758523347
transform 1 0 60474 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_11
timestamp 1758523347
transform 1 0 54146 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_12
timestamp 1758523347
transform 1 0 66802 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_13
timestamp 1758523347
transform 1 0 73130 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_14
timestamp 1758523347
transform 1 0 79458 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_15
timestamp 1758523347
transform 1 0 85786 0 1 13737
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_16
timestamp 1758523347
transform 1 0 85786 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_17
timestamp 1758523347
transform 1 0 79458 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_18
timestamp 1758523347
transform 1 0 79458 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_19
timestamp 1758523347
transform 1 0 85786 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_20
timestamp 1758523347
transform 1 0 73130 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_21
timestamp 1758523347
transform 1 0 73130 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_22
timestamp 1758523347
transform 1 0 66802 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_23
timestamp 1758523347
transform 1 0 66802 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_24
timestamp 1758523347
transform 1 0 60474 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_25
timestamp 1758523347
transform 1 0 60474 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_26
timestamp 1758523347
transform 1 0 54146 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_27
timestamp 1758523347
transform 1 0 54146 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_28
timestamp 1758523347
transform 1 0 47818 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_29
timestamp 1758523347
transform 1 0 41490 0 1 20905
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_30
timestamp 1758523347
transform 1 0 41490 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_31
timestamp 1758523347
transform 1 0 47818 0 1 24489
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_32
timestamp 1758523347
transform 1 0 41490 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_33
timestamp 1758523347
transform 1 0 41490 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_34
timestamp 1758523347
transform 1 0 47818 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_35
timestamp 1758523347
transform 1 0 54146 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_36
timestamp 1758523347
transform 1 0 54146 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_37
timestamp 1758523347
transform 1 0 47818 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_38
timestamp 1758523347
transform 1 0 60474 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_39
timestamp 1758523347
transform 1 0 60474 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_40
timestamp 1758523347
transform 1 0 66802 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_41
timestamp 1758523347
transform 1 0 73130 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_42
timestamp 1758523347
transform 1 0 73130 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_43
timestamp 1758523347
transform 1 0 66802 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_44
timestamp 1758523347
transform 1 0 79458 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_45
timestamp 1758523347
transform 1 0 79458 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_46
timestamp 1758523347
transform 1 0 85786 0 1 31657
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_47
timestamp 1758523347
transform 1 0 85786 0 1 28073
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_49
timestamp 1758523347
transform 1 0 85786 0 1 35241
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_50
timestamp 1758523347
transform 1 0 79458 0 1 38825
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_51
timestamp 1758523347
transform 1 0 79458 0 1 35241
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_52
timestamp 1758523347
transform 1 0 66802 0 1 38825
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_53
timestamp 1758523347
transform 1 0 66802 0 1 35241
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_54
timestamp 1758523347
transform 1 0 73130 0 1 38825
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_55
timestamp 1758523347
transform 1 0 73130 0 1 35241
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_56
timestamp 1758523347
transform 1 0 60474 0 1 38825
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_57
timestamp 1758523347
transform 1 0 60474 0 1 35241
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_58
timestamp 1758523347
transform 1 0 47818 0 1 38825
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_59
timestamp 1758523347
transform 1 0 47818 0 1 35241
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_60
timestamp 1758523347
transform 1 0 54146 0 1 38825
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_61
timestamp 1758523347
transform 1 0 54146 0 1 35241
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_62
timestamp 1758523347
transform 1 0 41490 0 1 38825
box -1114 -857 6338 3284
use unit_cell_aray  unit_cell_aray_63
timestamp 1758523347
transform 1 0 41490 0 1 35241
box -1114 -857 6338 3284
<< labels >>
flabel metal2 40544 16408 40824 16632 1 FreeSans 8000 0 0 0 D1
port 1 n
flabel metal2 40544 19992 40824 20216 1 FreeSans 8000 0 0 0 D2
port 2 n
flabel metal2 40544 23576 40824 23800 1 FreeSans 8000 0 0 0 D3
port 3 n
flabel metal2 40544 27160 40824 27384 1 FreeSans 8000 0 0 0 D4
port 4 n
flabel metal2 40544 30744 40824 30968 1 FreeSans 8000 0 0 0 D5
port 5 n
flabel metal2 40544 34328 40824 34552 1 FreeSans 8000 0 0 0 D6
port 6 n
flabel metal2 40544 37912 40824 38136 1 FreeSans 8000 0 0 0 D7
port 7 n
flabel metal2 40900 41730 41040 41990 1 FreeSans 8000 0 0 0 C1
port 8 n
flabel metal2 47230 41730 47370 41990 1 FreeSans 8000 0 0 0 C2
port 9 n
flabel metal2 53550 41730 53690 41990 1 FreeSans 8000 0 0 0 C3
port 10 n
flabel metal2 59880 41730 60020 41990 1 FreeSans 8000 0 0 0 C4
port 11 n
flabel metal2 66210 41730 66350 41990 1 FreeSans 8000 0 0 0 C5
port 12 n
flabel metal2 72530 41730 72670 41990 1 FreeSans 8000 0 0 0 C6
port 13 n
flabel metal2 78860 41730 79000 41990 1 FreeSans 8000 0 0 0 C7
port 14 n
flabel metal1 40210 40214 40421 40676 1 FreeSans 8000 0 0 0 CLK
port 15 n
flabel metal1 91723 41557 91934 42019 1 FreeSans 8000 0 0 0 OUTP
port 16 n
flabel metal1 92160 40164 92371 40626 1 FreeSans 8000 0 0 0 OUTN
port 17 n
flabel metal1 92631 38873 92842 39335 1 FreeSans 8000 0 0 0 VBIAS
port 18 n
flabel metal1 40829 12836 41513 13028 1 FreeSans 8000 0 0 0 VDD
port 19 n
flabel metal1 43470 41508 44154 41700 1 FreeSans 8000 0 0 0 VSS
port 20 n
<< end >>
