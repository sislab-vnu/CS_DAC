magic
tech gf180mcuD
magscale 1 10
timestamp 1754559251
<< pwell >>
rect -376 -185 1183 488
<< nmos >>
rect -238 240 -182 284
rect -14 240 42 284
rect 290 240 346 284
rect 466 240 522 284
rect 770 240 826 284
rect 994 240 1050 284
rect -238 0 -182 90
rect 0 0 360 90
rect 452 0 812 90
rect 994 0 1050 90
<< ndiff >>
rect 62 285 134 298
rect 62 284 75 285
rect -322 240 -238 284
rect -182 240 -136 284
rect -80 240 -14 284
rect 42 240 75 284
rect -80 90 -34 240
rect 62 239 75 240
rect 121 239 134 285
rect 62 226 134 239
rect 190 285 270 302
rect 190 239 207 285
rect 253 284 270 285
rect 366 287 446 304
rect 366 284 383 287
rect 253 240 290 284
rect 346 241 383 284
rect 429 284 446 287
rect 542 285 622 302
rect 542 284 559 285
rect 429 241 466 284
rect 346 240 466 241
rect 522 240 559 284
rect 253 239 270 240
rect 190 222 270 239
rect 366 224 446 240
rect 542 239 559 240
rect 605 239 622 285
rect 542 222 622 239
rect 678 285 750 298
rect 678 239 691 285
rect 737 284 750 285
rect 737 240 770 284
rect 826 240 892 284
rect 948 240 994 284
rect 1050 240 1134 284
rect 737 239 750 240
rect 678 226 750 239
rect 846 90 892 240
rect -284 0 -238 90
rect -182 0 -136 90
rect -80 0 0 90
rect 360 0 452 90
rect 812 0 892 90
rect 948 0 994 90
rect 1050 0 1096 90
rect 384 -56 428 0
rect 380 -66 432 -56
rect 366 -79 446 -66
rect 366 -125 383 -79
rect 429 -125 446 -79
rect 366 -138 446 -125
<< ndiffc >>
rect 75 239 121 285
rect 207 239 253 285
rect 383 241 429 287
rect 559 239 605 285
rect 691 239 737 285
rect 383 -125 429 -79
<< polysilicon >>
rect -26 407 54 424
rect -26 361 -9 407
rect 37 361 54 407
rect -26 344 54 361
rect 278 407 358 424
rect 278 361 295 407
rect 341 361 358 407
rect 278 344 358 361
rect 454 407 534 424
rect 454 361 471 407
rect 517 361 534 407
rect 454 344 534 361
rect 758 407 838 424
rect 758 361 775 407
rect 821 361 838 407
rect 758 344 838 361
rect -238 284 -182 328
rect -14 284 42 344
rect -238 90 -182 240
rect -14 194 42 240
rect 290 284 346 344
rect 466 284 522 344
rect 290 194 346 240
rect 466 194 522 240
rect 770 284 826 344
rect 994 284 1050 328
rect 770 194 826 240
rect 0 136 42 194
rect 324 136 488 146
rect 770 136 812 194
rect 0 110 812 136
rect 0 90 360 110
rect 452 90 812 110
rect 994 90 1050 240
rect -238 -46 -182 0
rect 0 -46 360 0
rect -246 -58 -174 -46
rect 452 -46 812 0
rect 994 -46 1050 0
rect -246 -104 -233 -58
rect -187 -104 -174 -58
rect 986 -58 1058 -46
rect -246 -118 -174 -104
rect 986 -104 999 -58
rect 1045 -104 1058 -58
rect 986 -118 1058 -104
<< polycontact >>
rect -9 361 37 407
rect 295 361 341 407
rect 471 361 517 407
rect 775 361 821 407
rect -233 -104 -187 -58
rect 999 -104 1045 -58
<< metal1 >>
rect -24 407 52 422
rect -24 361 -9 407
rect 37 361 52 407
rect -24 346 52 361
rect 280 407 356 422
rect 280 361 295 407
rect 341 361 356 407
rect 280 346 356 361
rect 456 407 532 422
rect 456 361 471 407
rect 517 361 532 407
rect 456 346 532 361
rect 760 407 836 422
rect 760 361 775 407
rect 821 361 836 407
rect 760 346 836 361
rect 75 285 121 296
rect 75 168 121 239
rect 192 285 268 300
rect 192 239 207 285
rect 253 239 268 285
rect 192 224 268 239
rect 383 287 429 298
rect 383 168 429 241
rect 544 285 620 300
rect 544 239 559 285
rect 605 239 620 285
rect 544 224 620 239
rect 691 285 737 296
rect 691 168 737 239
rect 75 122 737 168
rect -272 -58 1082 -24
rect -272 -104 -233 -58
rect -187 -79 999 -58
rect -187 -104 383 -79
rect -272 -125 383 -104
rect 429 -104 999 -79
rect 1045 -104 1082 -58
rect 429 -125 1082 -104
rect -272 -144 1082 -125
<< labels >>
flabel metal1 280 346 356 422 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 456 346 532 422 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 192 224 268 300 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 544 224 620 300 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 760 346 836 422 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 -24 346 52 422 1 FreeSans 400 0 0 0 VBIAS
port 6 nsew power bidirectional
flabel metal1 -187 -79 999 -24 1 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional
flabel pwell 841 -146 971 -20 1 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
<< end >>
