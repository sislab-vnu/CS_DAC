magic
tech gf180mcuD
magscale 1 10
timestamp 1754638763
<< isosubstrate >>
rect -416 1458 825 1490
rect -416 1439 94 1458
rect 170 1439 238 1458
rect 314 1439 825 1458
rect -416 820 825 1439
<< pwell >>
rect -416 1458 825 1490
rect -416 1439 94 1458
rect 170 1439 238 1458
rect 314 1439 825 1458
rect -416 820 825 1439
<< nmos >>
rect -294 1214 -234 1334
rect 102 1214 162 1334
rect 246 1214 306 1334
rect 642 1214 702 1334
rect -294 1002 -234 1064
rect -40 1002 20 1064
rect 106 1004 162 1060
rect 246 1004 302 1060
rect 386 1002 446 1064
rect 642 1002 702 1064
<< ndiff >>
rect -340 1214 -294 1334
rect -234 1214 -188 1334
rect 10 1317 102 1334
rect 10 1271 27 1317
rect 73 1271 102 1317
rect 10 1254 102 1271
rect 56 1214 102 1254
rect 162 1214 246 1334
rect 306 1317 398 1334
rect 306 1271 335 1317
rect 381 1271 398 1317
rect 306 1254 398 1271
rect 306 1214 352 1254
rect 596 1214 642 1334
rect 702 1214 748 1334
rect -132 1064 -60 1074
rect -340 1002 -294 1064
rect -234 1002 -188 1064
rect -132 1061 -40 1064
rect -132 1015 -119 1061
rect -73 1015 -40 1061
rect -132 1002 -40 1015
rect 20 1060 70 1064
rect 182 1060 226 1214
rect 468 1064 540 1074
rect 338 1060 386 1064
rect 20 1004 106 1060
rect 162 1004 246 1060
rect 302 1004 386 1060
rect 20 1002 86 1004
rect 42 928 86 1002
rect 322 1002 386 1004
rect 446 1061 540 1064
rect 446 1015 481 1061
rect 527 1015 540 1061
rect 446 1002 540 1015
rect 596 1002 642 1064
rect 702 1002 748 1064
rect 322 928 366 1002
rect 42 884 366 928
<< ndiffc >>
rect 27 1271 73 1317
rect 335 1271 381 1317
rect -119 1015 -73 1061
rect 481 1015 527 1061
<< polysilicon >>
rect 92 1443 172 1460
rect 92 1397 109 1443
rect 155 1397 172 1443
rect 92 1380 172 1397
rect 236 1443 316 1460
rect 236 1397 253 1443
rect 299 1397 316 1443
rect 236 1380 316 1397
rect -294 1334 -234 1380
rect 102 1334 162 1380
rect 246 1334 306 1380
rect 642 1334 702 1380
rect -294 1064 -234 1214
rect -118 1179 -38 1196
rect -118 1133 -101 1179
rect -55 1152 -38 1179
rect 102 1168 162 1214
rect -55 1133 -4 1152
rect -118 1120 -4 1133
rect -118 1116 162 1120
rect -40 1084 162 1116
rect -40 1064 20 1084
rect 106 1060 162 1084
rect 246 1168 306 1214
rect 446 1179 526 1196
rect 446 1152 463 1179
rect 410 1133 463 1152
rect 509 1133 526 1179
rect 410 1120 526 1133
rect 246 1116 526 1120
rect 246 1084 446 1116
rect 246 1060 302 1084
rect 386 1064 446 1084
rect 642 1064 702 1214
rect -294 958 -234 1002
rect -300 945 -228 958
rect -40 956 20 1002
rect -300 899 -287 945
rect -241 899 -228 945
rect -300 886 -228 899
rect 106 984 162 1004
rect 246 984 302 1004
rect 106 948 302 984
rect 386 956 446 1002
rect 642 956 702 1002
rect 636 943 708 956
rect 636 897 649 943
rect 695 897 708 943
rect 636 884 708 897
<< polycontact >>
rect 109 1397 155 1443
rect 253 1397 299 1443
rect -101 1133 -55 1179
rect 463 1133 509 1179
rect -287 899 -241 945
rect 649 897 695 943
<< metal1 >>
rect 94 1443 170 1458
rect 94 1397 109 1443
rect 155 1397 170 1443
rect 94 1382 170 1397
rect 238 1443 314 1458
rect 238 1397 253 1443
rect 299 1397 314 1443
rect 238 1382 314 1397
rect 12 1317 88 1332
rect 12 1271 27 1317
rect 73 1271 88 1317
rect 12 1256 88 1271
rect 320 1317 396 1332
rect 320 1271 335 1317
rect 381 1271 396 1317
rect 320 1256 396 1271
rect -116 1179 -40 1194
rect -116 1133 -101 1179
rect -55 1133 -40 1179
rect -116 1118 -40 1133
rect 448 1179 524 1194
rect 448 1133 463 1179
rect 509 1133 524 1179
rect 448 1118 524 1133
rect -119 1061 -73 1072
rect -119 980 -73 1015
rect 481 1061 527 1072
rect 481 980 527 1015
rect -340 945 758 980
rect -340 899 -287 945
rect -241 943 758 945
rect -241 899 649 943
rect -340 897 649 899
rect 695 897 758 943
rect -340 860 758 897
<< labels >>
flabel metal1 -116 1118 -40 1194 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 448 1118 524 1194 1 FreeSans 400 0 0 0 VBIAS
port 6 nsew power bidirectional
flabel metal1 -146 860 547 980 1 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional
flabel pwell 502 844 581 990 1 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
flabel metal1 94 1382 170 1458 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 238 1382 314 1458 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 12 1256 88 1332 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 320 1256 396 1332 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
<< end >>
