magic
tech gf180mcuD
magscale 1 10
timestamp 1756615742
<< nwell >>
rect 1741 4648 1915 4704
rect 1338 3800 1414 3876
<< psubdiff >>
rect 1957 5208 2057 5232
rect 1957 5152 1978 5208
rect 2034 5152 2057 5208
rect 1957 5132 2057 5152
rect 2016 3417 2116 3440
rect 2016 3360 2041 3417
rect 2097 3360 2116 3417
rect 2016 3340 2116 3360
rect 1937 1624 2037 1648
rect 1937 1568 1960 1624
rect 2016 1568 2037 1624
rect 1937 1548 2037 1568
rect 2009 -171 2109 -144
rect 2009 -227 2034 -171
rect 2090 -227 2109 -171
rect 2009 -244 2109 -227
<< nsubdiff >>
rect 1956 5993 2056 6016
rect 1956 5937 1983 5993
rect 2039 5937 2056 5993
rect 1956 5916 2056 5937
rect 2000 4200 2100 4224
rect 2000 4144 2019 4200
rect 2075 4144 2100 4200
rect 2000 4124 2100 4144
rect 1960 2408 2060 2432
rect 1960 2352 1981 2408
rect 2037 2352 2060 2408
rect 1960 2332 2060 2352
rect 2016 616 2116 640
rect 2016 560 2040 616
rect 2096 560 2116 616
rect 2016 540 2116 560
<< psubdiffcont >>
rect 1978 5152 2034 5208
rect 2041 3360 2097 3417
rect 1960 1568 2016 1624
rect 2034 -227 2090 -171
<< nsubdiffcont >>
rect 1983 5937 2039 5993
rect 2019 4144 2075 4200
rect 1981 2352 2037 2408
rect 2040 560 2096 616
<< metal1 >>
rect 336 5488 504 6384
rect 3528 6160 3696 6384
rect 2340 6104 2352 6160
rect 2408 6104 3696 6160
rect 1681 5544 2150 5600
rect 336 5432 1176 5488
rect 336 4704 504 5432
rect 336 4648 1176 4704
rect 336 3696 504 4648
rect 3528 4480 3696 6104
rect 3528 4424 3584 4480
rect 3640 4424 3696 4480
rect 3528 4368 3696 4424
rect 2408 4364 3696 4368
rect 2408 4312 2466 4364
rect 2518 4312 3696 4364
rect 1700 3752 2278 3808
rect 336 3640 1165 3696
rect 336 1904 504 3640
rect 3528 3136 3696 4312
rect 3528 3080 3584 3136
rect 3640 3080 3696 3136
rect 3528 2576 3696 3080
rect 2340 2520 2352 2576
rect 2408 2520 3696 2576
rect 1680 1904 2173 1960
rect 336 1848 1173 1904
rect 336 112 504 1848
rect 716 896 728 952
rect 784 896 2464 952
rect 2520 896 2532 952
rect 3528 784 3696 2520
rect 1332 728 1344 784
rect 1400 728 3696 784
rect 1729 112 2016 168
rect 2072 112 2279 168
rect 336 56 1164 112
rect 336 -337 504 56
rect 3528 -337 3696 728
<< via1 >>
rect 2352 6104 2408 6160
rect 1512 5936 1624 5992
rect 2352 5768 2408 5824
rect 1344 5600 1400 5656
rect 2688 5544 2744 5600
rect 2520 5152 2632 5208
rect 1686 4648 1742 4704
rect 1344 4424 1400 4480
rect 3584 4424 3640 4480
rect 2466 4312 2518 4364
rect 1512 4200 1624 4256
rect 2464 3976 2520 4032
rect 1344 3808 1400 3864
rect 2800 3752 2856 3808
rect 2520 3360 2632 3416
rect 1126 3080 1182 3136
rect 3584 3080 3640 3136
rect 1680 2912 1736 2968
rect 2352 2520 2408 2576
rect 1512 2408 1624 2464
rect 2352 2184 2408 2240
rect 1344 2016 1400 2072
rect 2688 1960 2744 2016
rect 2520 1568 2632 1624
rect 728 896 784 952
rect 2464 896 2520 952
rect 1344 728 1400 784
rect 1512 560 1624 616
rect 1344 392 1400 448
rect 2464 395 2520 451
rect 2016 112 2072 168
rect 2806 141 2862 197
rect 2520 -224 2632 -168
<< metal2 >>
rect 672 5656 840 6384
rect 2340 6160 2416 6170
rect 2340 6104 2352 6160
rect 2408 6104 2416 6160
rect 2340 6094 2416 6104
rect 1501 5992 1632 6002
rect 1501 5936 1512 5992
rect 1624 5936 1632 5992
rect 1501 5928 1632 5936
rect 2352 5834 2408 6094
rect 2344 5824 2420 5834
rect 2344 5768 2352 5824
rect 2408 5768 2420 5824
rect 2344 5758 2420 5768
rect 1336 5656 1412 5667
rect 672 5600 1344 5656
rect 1400 5600 1412 5656
rect 672 3864 840 5600
rect 1336 5591 1412 5600
rect 2678 5600 2754 5611
rect 2678 5544 2688 5600
rect 2744 5544 3920 5600
rect 2678 5535 2754 5544
rect 2508 5208 2644 5215
rect 2508 5152 2520 5208
rect 2632 5152 2644 5208
rect 2508 5143 2644 5152
rect 1677 4704 1753 4715
rect 1677 4648 1686 4704
rect 1742 4648 3920 4704
rect 1677 4639 1753 4648
rect 1336 4480 1412 4491
rect 3574 4480 3650 4491
rect 1336 4424 1344 4480
rect 1400 4424 3584 4480
rect 3640 4424 3650 4480
rect 1336 4415 1412 4424
rect 3574 4415 3650 4424
rect 2426 4364 2558 4368
rect 2426 4312 2466 4364
rect 2518 4312 2558 4364
rect 1503 4256 1632 4264
rect 1503 4200 1512 4256
rect 1624 4200 1632 4256
rect 1503 4189 1632 4200
rect 2464 4041 2520 4312
rect 2454 4032 2530 4041
rect 2454 3976 2464 4032
rect 2520 3976 2530 4032
rect 2454 3965 2530 3976
rect 1338 3864 1414 3876
rect 672 3808 1344 3864
rect 1400 3808 1414 3864
rect 672 2072 840 3808
rect 1338 3800 1414 3808
rect 2792 3808 2868 3819
rect 2792 3752 2800 3808
rect 2856 3752 3920 3808
rect 2792 3743 2868 3752
rect 2506 3416 2641 3424
rect 2506 3360 2520 3416
rect 2632 3360 2641 3416
rect 2506 3352 2641 3360
rect 1116 3136 1192 3147
rect 3573 3136 3649 3146
rect 1116 3080 1126 3136
rect 1182 3080 3584 3136
rect 3640 3080 3649 3136
rect 1116 3071 1192 3080
rect 3573 3070 3649 3080
rect 1671 2968 1747 2979
rect 1671 2912 1680 2968
rect 1736 2912 3920 2968
rect 1671 2903 1747 2912
rect 2340 2576 2416 2587
rect 2340 2520 2352 2576
rect 2408 2520 2416 2576
rect 2340 2511 2416 2520
rect 1503 2464 1632 2475
rect 1503 2408 1512 2464
rect 1624 2408 1632 2464
rect 1503 2400 1632 2408
rect 2352 2252 2408 2511
rect 2342 2240 2418 2252
rect 2342 2184 2352 2240
rect 2408 2184 2418 2240
rect 2342 2176 2418 2184
rect 1334 2072 1410 2084
rect 672 2016 1344 2072
rect 1400 2016 1410 2072
rect 672 952 840 2016
rect 1334 2008 1410 2016
rect 2680 2016 2756 2026
rect 2680 1960 2688 2016
rect 2744 1960 3920 2016
rect 2680 1950 2756 1960
rect 2512 1624 2641 1633
rect 2512 1568 2520 1624
rect 2632 1568 2641 1624
rect 2512 1559 2641 1568
rect 672 896 728 952
rect 784 896 840 952
rect 672 -337 840 896
rect 2016 1064 3920 1120
rect 1334 784 1410 794
rect 1334 728 1344 784
rect 1400 728 1410 784
rect 1334 718 1410 728
rect 1344 458 1400 718
rect 1501 616 1633 625
rect 1501 560 1512 616
rect 1624 560 1633 616
rect 1501 547 1633 560
rect 1334 448 1410 458
rect 1334 392 1344 448
rect 1400 392 1410 448
rect 1334 382 1410 392
rect 2016 178 2072 1064
rect 2453 952 2529 962
rect 2453 896 2464 952
rect 2520 896 2529 952
rect 2453 886 2529 896
rect 2464 461 2520 886
rect 2454 451 2530 461
rect 2454 395 2464 451
rect 2520 395 2530 451
rect 2454 385 2530 395
rect 2794 197 2874 210
rect 2005 168 2081 178
rect 2005 112 2016 168
rect 2072 112 2081 168
rect 2794 141 2806 197
rect 2862 141 3920 197
rect 2794 134 2874 141
rect 2005 102 2081 112
rect 2512 -168 2641 -160
rect 2512 -224 2520 -168
rect 2632 -224 2641 -168
rect 2512 -233 2641 -224
<< via2 >>
rect 1512 5936 1624 5992
rect 2520 5152 2632 5208
rect 1512 4200 1624 4256
rect 2520 3360 2632 3416
rect 1512 2408 1624 2464
rect 2520 1568 2632 1624
rect 1512 560 1624 616
rect 2520 -224 2632 -168
<< metal3 >>
rect 1456 5992 1680 6440
rect 1456 5936 1512 5992
rect 1624 5936 1680 5992
rect 1456 4256 1680 5936
rect 1456 4200 1512 4256
rect 1624 4200 1680 4256
rect 1456 2464 1680 4200
rect 1456 2408 1512 2464
rect 1624 2408 1680 2464
rect 1456 616 1680 2408
rect 1456 560 1512 616
rect 1624 560 1680 616
rect 1456 -336 1680 560
rect 2464 5208 2688 6440
rect 2464 5152 2520 5208
rect 2632 5152 2688 5208
rect 2464 3416 2688 5152
rect 2464 3360 2520 3416
rect 2632 3360 2688 3416
rect 2464 1624 2688 3360
rect 2464 1568 2520 1624
rect 2632 1568 2688 1624
rect 2464 -168 2688 1568
rect 2464 -224 2520 -168
rect 2632 -224 2688 -168
rect 2464 -336 2688 -224
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 982 0 1 5182
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_1
timestamp 1753044640
transform 1 0 982 0 -1 5070
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_2
timestamp 1753044640
transform 1 0 1990 0 1 5182
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_3
timestamp 1753044640
transform 1 0 982 0 1 1598
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_4
timestamp 1753044640
transform 1 0 2102 0 1 3390
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 982 0 -1 3278
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2102 0 1 -194
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_1
timestamp 1753044640
transform 1 0 982 0 1 3390
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_2
timestamp 1753044640
transform 1 0 1990 0 1 1598
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_4
timestamp 1753044640
transform 1 0 982 0 1 -194
box -86 -86 1206 870
<< labels >>
flabel metal2 672 6160 840 6384 1 FreeSans 3200 0 0 0 X0
port 1 n
flabel metal1 336 5152 504 5376 1 FreeSans 3200 0 0 0 X1
port 2 n
flabel metal2 3752 5544 3920 5600 1 FreeSans 3200 0 0 0 D7
port 10 n
flabel metal2 3752 4648 3920 4704 1 FreeSans 3200 0 0 0 D6
port 9 n
flabel metal2 3752 3752 3920 3808 1 FreeSans 3200 0 0 0 D5
port 8 n
flabel metal2 3752 2912 3920 2968 1 FreeSans 3200 0 0 0 D4
port 7 n
flabel metal2 3752 1960 3920 2016 1 FreeSans 3200 0 0 0 D3
port 6 n
flabel metal2 3752 1064 3920 1120 1 FreeSans 3200 0 0 0 D2
port 5 n
flabel metal1 3528 6160 3696 6384 1 FreeSans 3200 0 0 0 X2
port 3 n
flabel metal2 3752 141 3920 197 1 FreeSans 3200 0 0 0 D1
port 4 n
rlabel metal2 672 -337 840 6160 1 X0
port 1 n
rlabel metal1 336 5376 504 6384 1 X1
port 2 n
rlabel metal1 336 -337 504 5152 1 X1
port 2 n
rlabel metal1 3528 -337 3696 6160 1 X2
port 3 n
flabel metal3 1456 -336 1680 6440 1 FreeSans 3200 0 0 0 VDD
port 11 n
flabel metal3 2464 -336 2688 6440 1 FreeSans 3200 0 0 0 VSS
port 12 n
<< end >>
