** sch_path: /home/ducluong/CS_DAC/xschem/CS_Switch_1x.sch
.subckt CS_Switch_1x OUTN OUTP INP INN VBIAS VSS
*.PININFO INP:I INN:I OUTP:O OUTN:O VBIAS:B VSS:B
M1 net1 VBIAS net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 m=1
M2 OUTN INN net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 m=1
M3 net2 VBIAS VSS VSS nfet_03v3 L=2.2u W=0.22u nf=1 m=1
M4 OUTP INP net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 m=1
.ends
.end
