* NGSPICE file created from CS_Switch_16x2.ext - technology: gf180mcuD

.subckt CS_Switch_16x2 INP INN OUTP OUTN VBIAS VSS
X0 a_186_832# VBIAS a_64_826# VSS nfet_03v3 ad=0.1763p pd=1.32u as=99.299995f ps=0.95u w=0.56u l=0.28u
X1 a_64_826# VBIAS VSS VSS nfet_03v3 ad=99.299995f pd=0.95u as=0.1958p ps=1.6u w=0.62u l=0.3u
X2 a_334_832# VBIAS a_186_832# VSS nfet_03v3 ad=99.299995f pd=0.95u as=0.1763p ps=1.32u w=0.56u l=0.28u
X3 a_668_826# VSS VSS VSS nfet_03v3 ad=0.1426p pd=1.7u as=0.1958p ps=1.6u w=0.62u l=0.3u
X4 OUTN INN a_186_832# VSS nfet_03v3 ad=0.405p pd=1.95u as=0.23505p ps=1.76u w=0.6u l=0.3u
X5 VSS VBIAS a_334_832# VSS nfet_03v3 ad=0.1958p pd=1.6u as=99.299995f ps=0.95u w=0.62u l=0.3u
X6 a_668_1100# VSS OUTN VSS nfet_03v3 ad=0.138p pd=1.66u as=0.405p ps=1.95u w=0.6u l=0.3u
X7 VSS VSS a_n250_826# VSS nfet_03v3 ad=0.1958p pd=1.6u as=0.1426p ps=1.7u w=0.62u l=0.3u
X8 a_186_832# INP OUTP VSS nfet_03v3 ad=0.23505p pd=1.76u as=0.405p ps=1.95u w=0.6u l=0.3u
X9 OUTP VSS a_n250_1100# VSS nfet_03v3 ad=0.405p pd=1.95u as=0.138p ps=1.66u w=0.6u l=0.3u
C0 INP a_186_832# 5.25e-19
C1 a_186_832# VBIAS 0.002221f
C2 INP OUTN 0.001145f
C3 OUTN VBIAS 0.029999f
C4 INP INN 0.073624f
C5 INN VBIAS 0.020299f
C6 INP OUTP 0.002809f
C7 OUTP VBIAS 0.029999f
C8 OUTN a_668_1100# 0.001132f
C9 a_334_832# INN 2.43e-19
C10 OUTP a_n250_1100# 0.001132f
C11 INP VBIAS 0.020299f
C12 a_186_832# OUTN 0.002131f
C13 a_186_832# INN 5.25e-19
C14 a_186_832# OUTP 0.002131f
C15 OUTN INN 0.002809f
C16 OUTP OUTN 0.010625f
C17 INP a_64_826# 2.43e-19
C18 OUTP INN 0.001145f
C19 VBIAS VSS 0.771642f
C20 OUTN VSS 0.040088f
C21 OUTP VSS 0.040088f
C22 INN VSS 0.198651f
C23 INP VSS 0.198651f
C24 a_668_826# VSS 0.003029f
C25 a_334_832# VSS 0.004835f
C26 a_64_826# VSS 0.004835f
C27 a_n250_826# VSS 0.003029f
C28 a_668_1100# VSS 0.001094f
C29 a_186_832# VSS 0.010381f
C30 a_n250_1100# VSS 0.001094f
.ends

