** sch_path: /home/ducluong/CS_DAC/xschem/CS_DAC_10b.sch
**.subckt CS_DAC_10b
V1 vcc GND 3.3
V10 VBIAS GND 1.8
V2 X1 GND PULSE(0 3.3 0 1n 1n 4n 10n)
V5 X2 GND PULSE(0 3.3 0 1n 1n 9n 20n)
V6 X3 GND PULSE(0 3.3 0 1n 1n 19n 40n)
V7 X4 GND PULSE(0 3.3 0 1n 1n 39n 80n)
V8 X5 GND PULSE(0 3.3 0 1n 1n 79n 160n)
V9 X6 GND PULSE(0 3.3 0 1n 1n 159n 320n)
V11 X7 GND PULSE(0 3.3 0 1n 1n 319n 640n)
V12 X8 GND PULSE(0 3.3 0 1n 1n 639n 1280n)
V13 X9 GND PULSE(0 3.3 0 1n 1n 1279n 2560n)
V14 X10 GND PULSE(0 3.3 0 1n 1n 2559n 5120n)
V15 CLK GND PULSE(0 3.3 2n 1n 1n 4n 10n)
x1 X1 X2 X3 X4 net16 net15 VBIAS CLK vcc GND 4LSB_weighted_binary
x2 net14 net13 net12 net11 net10 net9 net8 net1 net2 net3 net4 net5 net6 net7 CLK net15 net16 VBIAS vcc GND 6MSB_matrix
x3 X8 X9 X10 net1 net3 net4 net5 net6 net2 net7 vcc GND thermometter_decoder
x4 X5 X6 X7 net14 net12 net11 net10 net9 net13 net8 vcc GND thermometter_decoder
R1 vcc net15 0 m=1
R2 vcc net16 0 m=1
**** begin user architecture code

.include /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.tech/ngspice/smbb000149.ngspice typical

 .include /home/ducluong/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/spice/gf180mcu_fd_sc_mcu7t5v0.spice


.save @R1[i] @R2[i] @R3[i] @R4[i]
.control
set wr_vecnames
set wr_singlescale
tran 1n 5120n
run
wrdata /home/ducluong/CS_DAC/spice/CS_DAC_10b.raw @R1[i] @R2[i]
.endc


**** end user architecture code
**.ends

* expanding   symbol:  4LSB_weighted_binary.sym # of pins=10
** sym_path: /home/ducluong/CS_DAC/xschem/4LSB_weighted_binary.sym
** sch_path: /home/ducluong/CS_DAC/xschem/4LSB_weighted_binary.sch
.subckt 4LSB_weighted_binary D1 D2 D3 D4 OUTP OUTN VBIAS CLK VDD VSS
*.ipin D1
*.ipin D2
*.ipin D3
*.ipin D4
*.opin OUTP
*.opin OUTN
*.opin VBIAS
*.ipin CLK
*.opin VDD
*.opin VSS
x5 D3 CLK net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
x6 D1 CLK net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
x7 D2 CLK net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
x8 D4 CLK net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
x9 net1 net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
x10 net2 net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
x11 net3 net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
x12 net4 net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
x1 net2 net6 OUTP OUTN VBIAS VSS CS_Switch_1x1
x2 net3 net7 OUTP OUTN VBIAS VSS CS_Switch_2x2
x3 net1 net5 OUTP OUTN VBIAS VSS CS_Switch_4x2
x4 net4 net8 OUTP OUTN VBIAS VSS CS_Switch_8x2
.ends


* expanding   symbol:  6MSB_matrix.sym # of pins=20
** sym_path: /home/ducluong/CS_DAC/xschem/6MSB_matrix.sym
** sch_path: /home/ducluong/CS_DAC/xschem/6MSB_matrix.sch
.subckt 6MSB_matrix C1 C2 C3 C4 C5 C6 C7 D1 D2 D3 D4 D5 D6 D7 CLK OUTP OUTN VBIAS VDD VSS
*.ipin D1
*.ipin D2
*.ipin D3
*.ipin D4
*.ipin D5
*.ipin D6
*.ipin D7
*.ipin C1
*.ipin C2
*.ipin C3
*.ipin C4
*.ipin C5
*.ipin C6
*.ipin C7
*.ipin CLK
*.iopin OUTP
*.iopin OUTN
*.iopin VBIAS
*.iopin VDD
*.iopin VSS
x7 C7 CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
x8 VSS CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
x9 C1 CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x10 C2 CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x11 C3 CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x12 C4 CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x13 C5 CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x14 C6 CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x15 C7 CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x16 VSS CLK OUTP OUTN VBIAS VDD D1 D2 VSS unit_cell_aray
x17 C1 CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x18 C2 CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x19 C3 CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x20 C4 CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x21 C5 CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x22 C6 CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x23 C7 CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x24 VSS CLK OUTP OUTN VBIAS VDD D2 D3 VSS unit_cell_aray
x25 C1 CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x26 C2 CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x27 C3 CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x28 C4 CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x29 C5 CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x30 C6 CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x31 C7 CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x32 VSS CLK OUTP OUTN VBIAS VDD D3 D4 VSS unit_cell_aray
x33 C1 CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x34 C2 CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x35 C3 CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x36 C4 CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x37 C5 CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x38 C6 CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x39 C7 CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x40 VSS CLK OUTP OUTN VBIAS VDD D4 D5 VSS unit_cell_aray
x41 C1 CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x42 C2 CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x43 C3 CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x44 C4 CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x45 C5 CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x46 C6 CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x47 C7 CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x48 VSS CLK OUTP OUTN VBIAS VDD D5 D6 VSS unit_cell_aray
x49 C1 CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x50 C2 CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x51 C3 CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x52 C4 CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x53 C5 CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x54 C6 CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x55 C7 CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x56 VSS CLK OUTP OUTN VBIAS VDD D6 D7 VSS unit_cell_aray
x57 C1 CLK OUTP OUTN VBIAS VDD D7 VSS VSS unit_cell_aray
x58 C2 CLK OUTP OUTN VBIAS VDD D7 VSS VSS unit_cell_aray
x59 C3 CLK OUTP OUTN VBIAS VDD D7 VSS VSS unit_cell_aray
x60 C4 CLK OUTP OUTN VBIAS VDD D7 VSS VSS unit_cell_aray
x61 C5 CLK OUTP OUTN VBIAS VDD D7 VSS VSS unit_cell_aray
x62 C6 CLK OUTP OUTN VBIAS VDD D7 VSS VSS unit_cell_aray
x63 C7 CLK OUTP OUTN VBIAS VDD D7 VSS VSS unit_cell_aray
x1 C1 CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
x2 C2 CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
x3 C3 CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
x4 C4 CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
x5 C5 CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
x6 C6 CLK OUTP OUTN VBIAS VDD VDD D1 VSS unit_cell_aray
.ends


* expanding   symbol:  thermometter_decoder.sym # of pins=12
** sym_path: /home/ducluong/CS_DAC/xschem/thermometter_decoder.sym
** sch_path: /home/ducluong/CS_DAC/xschem/thermometter_decoder.sch
.subckt thermometter_decoder X0 X1 X2 D1 D3 D4 D5 D6 D2 D7 VDD VSS
*.ipin X0
*.ipin X1
*.ipin X2
*.opin D1
*.opin D2
*.opin D3
*.opin D4
*.opin D5
*.opin D6
*.opin D7
*.iopin VDD
*.iopin VSS
x3 X1 X2 D6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
x4 X1 X0 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
x5 net2 X2 D5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
x6 X2 D4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
x7 X1 X0 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
x8 net3 X2 D3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
x9 X1 X2 D2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
x10 D2 X0 D1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
x1 X1 X0 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
x2 net1 X2 D7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_2
.ends


* expanding   symbol:  CS_Switch_1x1.sym # of pins=6
** sym_path: /home/ducluong/CS_DAC/xschem/CS_Switch_1x1.sym
** sch_path: /home/ducluong/CS_DAC/xschem/CS_Switch_1x1.sch
.subckt CS_Switch_1x1 INP INN OUTP OUTN VBIAS VSS
*.ipin INP
*.ipin INN
*.opin OUTP
*.opin OUTN
*.iopin VBIAS
*.iopin VSS
XM3 net1 VBIAS net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net2 VBIAS VSS VSS nfet_03v3 L=2.2u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 OUTN INN net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 net1 INP OUTP VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  CS_Switch_2x2.sym # of pins=6
** sym_path: /home/ducluong/CS_DAC/xschem/CS_Switch_2x2.sym
** sch_path: /home/ducluong/CS_DAC/xschem/CS_Switch_2x2.sch
.subckt CS_Switch_2x2 INP INN OUTP OUTN VBIAS VSS
*.ipin INP
*.ipin INN
*.opin OUTP
*.opin OUTN
*.iopin VBIAS
*.iopin VSS
XM1 net1 VBIAS net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 OUTN INN net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 OUTP INP net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net2 VBIAS VSS VSS nfet_03v3 L=1.8u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  CS_Switch_4x2.sym # of pins=6
** sym_path: /home/ducluong/CS_DAC/xschem/CS_Switch_4x2.sym
** sch_path: /home/ducluong/CS_DAC/xschem/CS_Switch_4x2.sch
.subckt CS_Switch_4x2 INP INN OUTP OUTN VBIAS VSS
*.ipin INP
*.ipin INN
*.opin OUTP
*.opin OUTN
*.iopin VBIAS
*.iopin VSS
XM2 OUTP INP net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net1 VBIAS net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net2 VBIAS VSS VSS nfet_03v3 L=1.8u W=0.45u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net1 VBIAS net3 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 net1 INN OUTN VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM10 net3 VBIAS VSS VSS nfet_03v3 L=1.8u W=0.45u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  CS_Switch_8x2.sym # of pins=6
** sym_path: /home/ducluong/CS_DAC/xschem/CS_Switch_8x2.sym
** sch_path: /home/ducluong/CS_DAC/xschem/CS_Switch_8x2.sch
.subckt CS_Switch_8x2 INP INN OUTP OUTN VBIAS VSS
*.ipin INP
*.ipin INN
*.opin OUTP
*.opin OUTN
*.iopin VBIAS
*.iopin VSS
XM5 net1 VBIAS net2 VSS nfet_03v3 L=0.28u W=0.56u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net2 VBIAS VSS VSS nfet_03v3 L=0.3u W=0.62u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM1 OUTP INP net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 OUTN INN net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  unit_cell_aray.sym # of pins=9
** sym_path: /home/ducluong/CS_DAC/xschem/unit_cell_aray.sym
** sch_path: /home/ducluong/CS_DAC/xschem/unit_cell_aray.sch
.subckt unit_cell_aray Ci CLK OUTP OUTN VBIAS VDD Ri-1 Ri VSS
*.ipin Ci
*.ipin CLK
*.opin OUTP
*.opin OUTN
*.iopin VBIAS
*.iopin VDD
*.ipin Ri-1
*.ipin Ri
*.iopin VSS
x4 net1 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
x1 net3 CLK net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
x2 Ri Ci net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__or2_2
x3 net4 Ri-1 net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_2
x5 net1 net2 OUTP OUTN VBIAS VSS CS_Switch_16x2
.ends


* expanding   symbol:  CS_Switch_16x2.sym # of pins=6
** sym_path: /home/ducluong/CS_DAC/xschem/CS_Switch_16x2.sym
** sch_path: /home/ducluong/CS_DAC/xschem/CS_Switch_16x2.sch
.subckt CS_Switch_16x2 INP INN OUTP OUTN VBIAS VSS
*.ipin INP
*.ipin INN
*.opin OUTP
*.opin OUTN
*.iopin VBIAS
*.iopin VSS
XM2 net2 VBIAS VSS VSS nfet_03v3 L=0.3u W=0.62u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM1 net1 VBIAS net2 VSS nfet_03v3 L=0.28u W=0.56u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net1 VBIAS net3 VSS nfet_03v3 L=0.28u W=0.56u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 OUTN INN net1 VSS nfet_03v3 L=0.3u W=0.6u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net3 VBIAS VSS VSS nfet_03v3 L=0.3u W=0.62u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM9 OUTP INP net1 VSS nfet_03v3 L=0.3u W=0.6u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
