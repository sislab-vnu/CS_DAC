magic
tech gf180mcuD
magscale 1 10
timestamp 1758278152
<< isosubstrate >>
rect 8750 1010 8764 1152
rect 9350 966 9406 1130
rect 8735 504 8819 942
<< pwell >>
rect 8750 1010 8764 1152
rect 9350 966 9406 1130
rect 8735 504 8819 942
rect 8970 -113 9026 44
rect 9072 -125 9100 -81
rect 8744 -456 8763 -178
rect 8970 -216 9026 -187
rect 6805 -590 6870 -456
rect 8728 -590 9824 -456
rect 8744 -616 8763 -590
rect 10090 -1176 10146 -1120
rect 8741 -1575 8770 -1298
rect 6804 -1710 6870 -1575
rect 8728 -1710 10070 -1575
rect 8741 -1736 8770 -1710
rect 8750 -2344 8822 -2161
rect 8750 -2407 8954 -2344
rect 9343 -2378 9399 -2184
rect 8751 -2418 8954 -2407
rect 8729 -2603 8954 -2418
rect 8729 -2626 8826 -2603
rect 8748 -2649 8826 -2626
rect 6805 -2830 6870 -2649
rect 8728 -2830 10183 -2649
rect 8748 -2856 8826 -2830
<< psubdiff >>
rect 2672 623 2772 640
rect 2672 557 2691 623
rect 2751 557 2772 623
rect 2672 540 2772 557
rect 9530 537 9638 626
rect 2672 -503 2772 -480
rect 2672 -560 2692 -503
rect 2748 -560 2772 -503
rect 2672 -580 2772 -560
rect 9527 -589 9644 -485
rect 2672 -1622 2772 -1600
rect 2672 -1682 2694 -1622
rect 2753 -1682 2772 -1622
rect 2672 -1700 2772 -1682
rect 2672 -2736 2772 -2720
rect 2672 -2800 2689 -2736
rect 2750 -2800 2772 -2736
rect 2672 -2820 2772 -2800
<< nsubdiff >>
rect 2672 1407 2772 1424
rect 2672 1341 2690 1407
rect 2750 1341 2772 1407
rect 2672 1324 2772 1341
rect 2672 280 2772 304
rect 2672 223 2693 280
rect 2749 223 2772 280
rect 2672 204 2772 223
rect 2672 -840 2772 -816
rect 2672 -900 2691 -840
rect 2750 -900 2772 -840
rect 2672 -916 2772 -900
rect 2672 -1956 2772 -1936
rect 2672 -2020 2691 -1956
rect 2752 -2020 2772 -1956
rect 2672 -2036 2772 -2020
<< psubdiffcont >>
rect 2691 557 2751 623
rect 2692 -560 2748 -503
rect 2694 -1682 2753 -1622
rect 2689 -2800 2750 -2736
<< nsubdiffcont >>
rect 2690 1341 2750 1407
rect 2693 223 2749 280
rect 2691 -900 2750 -840
rect 2691 -2020 2752 -1956
<< metal1 >>
rect 2240 1020 2576 1680
rect 6777 1412 6899 1434
rect 5432 1344 5544 1400
rect 6836 1332 6899 1412
rect 6777 1314 6899 1332
rect 8943 1400 10072 1456
rect 10128 1400 10146 1456
rect 7907 1020 8096 1022
rect 2240 944 2801 1020
rect 5939 1008 6269 1014
rect 5936 952 6273 1008
rect 2240 -100 2576 944
rect 5939 931 6269 952
rect 8943 882 8999 1400
rect 10248 1288 10584 1624
rect 9350 1232 10584 1288
rect 9350 882 9406 1232
rect 9526 1064 10078 1120
rect 10134 1064 10146 1120
rect 8661 682 8741 683
rect 6806 530 6870 650
rect 8661 530 9781 682
rect 6800 301 6884 314
rect 5432 224 5544 280
rect 6822 221 6884 301
rect 6800 194 6884 221
rect 8970 280 10069 336
rect 10125 280 10146 336
rect 2240 -176 2803 -100
rect 5936 -139 6324 -112
rect 5944 -168 6260 -139
rect 2240 -1220 2576 -176
rect 8970 -216 9026 280
rect 10248 168 10584 1232
rect 9374 112 10584 168
rect 9374 -216 9430 112
rect 9552 -56 10078 0
rect 10134 -56 10146 0
rect 8728 -470 9824 -456
rect 6805 -590 6870 -470
rect 8657 -590 9824 -470
rect 6800 -823 6888 -806
rect 5432 -896 5544 -840
rect 6826 -903 6888 -823
rect 6800 -926 6888 -903
rect 9225 -840 10074 -784
rect 10130 -840 10146 -784
rect 2240 -1296 2802 -1220
rect 5929 -1288 6277 -1232
rect 2240 -2340 2576 -1296
rect 9225 -1327 9281 -840
rect 10248 -952 10584 112
rect 9642 -1008 10584 -952
rect 9642 -1327 9698 -1008
rect 9814 -1176 10076 -1120
rect 10132 -1176 10146 -1120
rect 8728 -1590 10070 -1575
rect 6804 -1710 6870 -1590
rect 8652 -1710 10070 -1590
rect 6799 -1947 6883 -1926
rect 5432 -2016 5544 -1960
rect 6830 -2027 6883 -1947
rect 6799 -2046 6883 -2027
rect 8970 -1960 10075 -1904
rect 10131 -1960 10146 -1904
rect 2240 -2352 2804 -2340
rect 2240 -2408 2806 -2352
rect 5936 -2407 6272 -2352
rect 2240 -2416 2804 -2408
rect 2240 -2968 2576 -2416
rect 8970 -2496 9026 -1960
rect 10248 -2072 10584 -1008
rect 9474 -2128 10584 -2072
rect 9474 -2496 9530 -2128
rect 9702 -2352 10133 -2296
rect 10189 -2352 10202 -2296
rect 8728 -2710 10183 -2649
rect 6805 -2830 6870 -2710
rect 8652 -2830 10183 -2710
rect 10248 -2912 10584 -2128
rect 10696 1456 11032 1624
rect 10696 1400 10808 1456
rect 10920 1400 11032 1456
rect 10696 336 11032 1400
rect 10696 280 10808 336
rect 10920 280 11032 336
rect 10696 -784 11032 280
rect 10696 -840 10808 -784
rect 10920 -840 11032 -784
rect 10696 -1904 11032 -840
rect 10696 -1960 10808 -1904
rect 10920 -1960 11032 -1904
rect 10696 -2912 11032 -1960
rect 11144 1120 11480 1624
rect 11144 1064 11256 1120
rect 11368 1064 11480 1120
rect 11144 0 11480 1064
rect 11144 -56 11256 0
rect 11368 -56 11480 0
rect 11144 -1120 11480 -56
rect 11144 -1176 11256 -1120
rect 11368 -1176 11480 -1120
rect 11144 -2296 11480 -1176
rect 11144 -2352 11256 -2296
rect 11368 -2352 11480 -2296
rect 11144 -2912 11480 -2352
<< via1 >>
rect 2838 1329 3000 1409
rect 4573 1333 4735 1413
rect 6674 1332 6836 1412
rect 10072 1400 10128 1456
rect 6397 1176 6453 1232
rect 8451 1057 8503 1109
rect 6496 952 6552 1008
rect 7018 924 7070 976
rect 7914 958 7966 1010
rect 3583 850 3639 906
rect 9064 1017 9120 1073
rect 9232 1017 9288 1073
rect 10078 1064 10134 1120
rect 7572 815 7624 867
rect 3768 549 3930 629
rect 5736 553 5898 633
rect 7744 549 7906 629
rect 2828 217 2990 297
rect 4600 213 4762 293
rect 6660 221 6822 301
rect 10069 280 10125 336
rect 6396 56 6452 112
rect 8459 -65 8511 -13
rect 6496 -179 6552 -123
rect 7021 -182 7073 -130
rect 7915 -166 7967 -114
rect 3582 -271 3638 -215
rect 9082 -84 9138 -28
rect 9258 -83 9314 -27
rect 10078 -56 10134 0
rect 7573 -298 7625 -246
rect 3772 -571 3934 -491
rect 5744 -567 5906 -487
rect 7752 -567 7914 -487
rect 2852 -903 3014 -823
rect 4584 -911 4746 -831
rect 6664 -903 6826 -823
rect 10074 -840 10130 -784
rect 6398 -1064 6454 -1008
rect 8457 -1182 8509 -1130
rect 6496 -1288 6552 -1232
rect 7021 -1295 7073 -1243
rect 7917 -1291 7969 -1239
rect 9345 -1195 9401 -1139
rect 9520 -1195 9576 -1139
rect 10076 -1176 10132 -1120
rect 3583 -1390 3639 -1334
rect 7573 -1416 7625 -1364
rect 3768 -1695 3930 -1615
rect 5728 -1687 5890 -1607
rect 7740 -1691 7902 -1611
rect 2836 -2023 2998 -1943
rect 4580 -2027 4742 -1947
rect 6668 -2027 6830 -1947
rect 10075 -1960 10131 -1904
rect 6395 -2240 6451 -2184
rect 8458 -2308 8510 -2256
rect 6496 -2408 6552 -2352
rect 7022 -2411 7074 -2359
rect 7917 -2409 7969 -2357
rect 3583 -2511 3639 -2455
rect 7573 -2538 7625 -2486
rect 9115 -2376 9171 -2320
rect 9343 -2378 9399 -2322
rect 10133 -2352 10189 -2296
rect 3764 -2810 3926 -2730
rect 5724 -2814 5886 -2734
rect 7752 -2810 7914 -2730
rect 10808 1400 10920 1456
rect 10808 280 10920 336
rect 10808 -840 10920 -784
rect 10808 -1960 10920 -1904
rect 11256 1064 11368 1120
rect 11256 -56 11368 0
rect 11256 -1176 11368 -1120
rect 11256 -2352 11368 -2296
<< metal2 >>
rect 10056 1456 10143 1467
rect 10780 1456 10947 1482
rect 2770 1409 3104 1434
rect 2770 1329 2838 1409
rect 3000 1329 3104 1409
rect 2770 1314 3104 1329
rect 4508 1413 4842 1434
rect 4508 1333 4573 1413
rect 4735 1333 4842 1413
rect 4508 1314 4842 1333
rect 6581 1412 6915 1434
rect 6581 1332 6674 1412
rect 6836 1332 6915 1412
rect 10056 1400 10072 1456
rect 10128 1400 10808 1456
rect 10920 1400 10976 1456
rect 10056 1384 10143 1400
rect 10780 1367 10947 1400
rect 6581 1314 6915 1332
rect 6387 1232 7981 1244
rect 6387 1176 6397 1232
rect 6453 1176 7981 1232
rect 6387 1161 7981 1176
rect 3576 906 3657 1132
rect 6478 1008 6564 1014
rect 7901 1010 7981 1161
rect 8436 1171 9298 1263
rect 8436 1109 8516 1171
rect 8436 1057 8451 1109
rect 8503 1057 8516 1109
rect 8436 1042 8516 1057
rect 9054 1073 9130 1082
rect 6478 952 6496 1008
rect 6552 976 7094 1008
rect 6552 952 7018 976
rect 6478 931 7018 952
rect 7011 924 7018 931
rect 7070 924 7094 976
rect 7901 958 7914 1010
rect 7966 958 7981 1010
rect 9054 1017 9064 1073
rect 9120 1017 9130 1073
rect 9054 1008 9130 1017
rect 7901 945 7981 958
rect 7011 912 7094 924
rect 3576 850 3583 906
rect 3639 850 3657 906
rect 9053 888 9130 1008
rect 9222 1073 9298 1171
rect 9222 1017 9232 1073
rect 9288 1017 9298 1073
rect 10063 1120 10146 1137
rect 11231 1120 11396 1147
rect 10063 1064 10078 1120
rect 10134 1064 11256 1120
rect 11368 1064 11424 1120
rect 10063 1048 10146 1064
rect 11231 1041 11396 1064
rect 9222 1006 9298 1017
rect 3576 832 3657 850
rect 7558 867 9130 888
rect 7558 815 7572 867
rect 7624 815 9130 867
rect 7558 803 9130 815
rect 3686 629 4020 650
rect 3686 549 3768 629
rect 3930 549 4020 629
rect 3686 530 4020 549
rect 5650 633 5984 650
rect 5650 553 5736 633
rect 5898 553 5984 633
rect 5650 530 5984 553
rect 7662 629 7996 650
rect 7662 549 7744 629
rect 7906 549 7996 629
rect 7662 530 7996 549
rect 10053 336 10136 355
rect 10778 336 10947 363
rect 2770 297 3104 314
rect 2770 217 2828 297
rect 2990 217 3104 297
rect 2770 194 3104 217
rect 4508 293 4842 314
rect 4508 213 4600 293
rect 4762 213 4842 293
rect 4508 194 4842 213
rect 6581 301 6915 314
rect 6581 221 6660 301
rect 6822 221 6915 301
rect 10053 280 10069 336
rect 10125 280 10808 336
rect 10920 280 10976 336
rect 10053 263 10136 280
rect 10778 250 10947 280
rect 6581 194 6915 221
rect 8446 124 8526 158
rect 6384 112 7979 122
rect 6384 56 6396 112
rect 6452 56 7979 112
rect 6384 46 7979 56
rect 3576 -215 3657 12
rect 7900 -96 7979 46
rect 8446 44 9325 124
rect 8446 -13 8526 44
rect 8446 -65 8459 -13
rect 8511 -65 8526 -13
rect 8446 -79 8526 -65
rect 9072 -28 9148 -18
rect 9072 -84 9082 -28
rect 9138 -84 9148 -28
rect 6481 -107 6564 -106
rect 6481 -123 7085 -107
rect 6481 -179 6496 -123
rect 6552 -130 7085 -123
rect 6552 -179 7021 -130
rect 6481 -182 7021 -179
rect 7073 -182 7085 -130
rect 7900 -114 7980 -96
rect 7900 -166 7915 -114
rect 7967 -166 7980 -114
rect 7900 -176 7980 -166
rect 6481 -189 7085 -182
rect 7005 -198 7085 -189
rect 3576 -271 3582 -215
rect 3638 -271 3657 -215
rect 9072 -237 9148 -84
rect 9248 -22 9325 44
rect 10061 0 10146 14
rect 11224 0 11393 27
rect 9248 -27 9324 -22
rect 9248 -83 9258 -27
rect 9314 -83 9324 -27
rect 10061 -56 10078 0
rect 10134 -56 11256 0
rect 11368 -56 11424 0
rect 10061 -69 10146 -56
rect 11224 -82 11393 -56
rect 9248 -94 9324 -83
rect 3576 -288 3657 -271
rect 7555 -246 9148 -237
rect 7555 -298 7573 -246
rect 7625 -298 9148 -246
rect 7555 -317 9148 -298
rect 3686 -491 4020 -470
rect 3686 -571 3772 -491
rect 3934 -571 4020 -491
rect 3686 -590 4020 -571
rect 5649 -487 5983 -470
rect 5649 -567 5744 -487
rect 5906 -567 5983 -487
rect 5649 -590 5983 -567
rect 7662 -487 7996 -470
rect 7662 -567 7752 -487
rect 7914 -567 7996 -487
rect 7662 -590 7996 -567
rect 10054 -784 10146 -761
rect 10778 -784 10950 -754
rect 2770 -823 3104 -806
rect 2770 -903 2852 -823
rect 3014 -903 3104 -823
rect 2770 -926 3104 -903
rect 4508 -831 4842 -806
rect 4508 -911 4584 -831
rect 4746 -911 4842 -831
rect 4508 -926 4842 -911
rect 6581 -823 6915 -806
rect 6581 -903 6664 -823
rect 6826 -903 6915 -823
rect 10054 -840 10074 -784
rect 10130 -840 10808 -784
rect 10920 -840 10976 -784
rect 10054 -861 10146 -840
rect 10778 -869 10950 -840
rect 6581 -926 6915 -903
rect 6387 -1008 7987 -993
rect 6387 -1064 6398 -1008
rect 6454 -1064 7987 -1008
rect 6387 -1073 7987 -1064
rect 3576 -1334 3657 -1108
rect 6482 -1230 7011 -1226
rect 6482 -1232 7091 -1230
rect 6482 -1288 6496 -1232
rect 6552 -1243 7091 -1232
rect 6552 -1288 7021 -1243
rect 6482 -1295 7021 -1288
rect 7073 -1295 7091 -1243
rect 6482 -1309 7091 -1295
rect 7907 -1239 7987 -1073
rect 8446 -1073 9591 -996
rect 8446 -1076 9274 -1073
rect 9466 -1076 9591 -1073
rect 8446 -1130 8526 -1076
rect 8446 -1182 8457 -1130
rect 8509 -1182 8526 -1130
rect 8446 -1196 8526 -1182
rect 9330 -1139 9410 -1129
rect 9330 -1195 9345 -1139
rect 9401 -1195 9410 -1139
rect 7907 -1291 7917 -1239
rect 7969 -1291 7987 -1239
rect 7907 -1300 7987 -1291
rect 6537 -1310 7091 -1309
rect 3576 -1390 3583 -1334
rect 3639 -1390 3657 -1334
rect 9330 -1357 9410 -1195
rect 9510 -1139 9591 -1076
rect 9510 -1195 9520 -1139
rect 9576 -1164 9591 -1139
rect 10064 -1120 10140 -1109
rect 11227 -1120 11399 -1090
rect 9576 -1195 9586 -1164
rect 10064 -1176 10076 -1120
rect 10132 -1176 11256 -1120
rect 11368 -1176 11424 -1120
rect 10064 -1185 10140 -1176
rect 9510 -1205 9586 -1195
rect 11227 -1207 11399 -1176
rect 3576 -1408 3657 -1390
rect 7560 -1364 9410 -1357
rect 7560 -1416 7573 -1364
rect 7625 -1416 9410 -1364
rect 7560 -1437 9410 -1416
rect 3686 -1615 4020 -1590
rect 3686 -1695 3768 -1615
rect 3930 -1695 4020 -1615
rect 3686 -1710 4020 -1695
rect 5649 -1607 5983 -1590
rect 5649 -1687 5728 -1607
rect 5890 -1687 5983 -1607
rect 5649 -1710 5983 -1687
rect 7662 -1611 7996 -1590
rect 7662 -1691 7740 -1611
rect 7902 -1691 7996 -1611
rect 7662 -1710 7996 -1691
rect 10059 -1904 10146 -1889
rect 10781 -1904 10944 -1881
rect 2770 -1943 3104 -1926
rect 2770 -2023 2836 -1943
rect 2998 -2023 3104 -1943
rect 2770 -2046 3104 -2023
rect 4508 -1947 4842 -1926
rect 4508 -2027 4580 -1947
rect 4742 -2027 4842 -1947
rect 4508 -2046 4842 -2027
rect 6581 -1947 6915 -1926
rect 6581 -2027 6668 -1947
rect 6830 -2027 6915 -1947
rect 10059 -1960 10075 -1904
rect 10131 -1960 10808 -1904
rect 10920 -1960 10976 -1904
rect 10059 -1974 10146 -1960
rect 10781 -1987 10944 -1960
rect 6581 -2046 6915 -2027
rect 8446 -2163 8526 -2162
rect 6383 -2184 7986 -2172
rect 3576 -2455 3657 -2228
rect 6383 -2240 6395 -2184
rect 6451 -2240 7986 -2184
rect 6383 -2252 7986 -2240
rect 6483 -2347 6564 -2346
rect 6483 -2352 7091 -2347
rect 6483 -2408 6496 -2352
rect 6552 -2359 7091 -2352
rect 6552 -2408 7022 -2359
rect 6483 -2411 7022 -2408
rect 7074 -2411 7091 -2359
rect 6483 -2427 7091 -2411
rect 7906 -2357 7986 -2252
rect 8446 -2242 9399 -2163
rect 8446 -2256 8526 -2242
rect 8446 -2308 8458 -2256
rect 8510 -2308 8526 -2256
rect 8446 -2328 8526 -2308
rect 9343 -2312 9399 -2242
rect 10122 -2296 10198 -2286
rect 11227 -2296 11396 -2268
rect 9105 -2320 9181 -2312
rect 7906 -2409 7917 -2357
rect 7969 -2409 7986 -2357
rect 7906 -2418 7986 -2409
rect 9105 -2376 9115 -2320
rect 9171 -2376 9181 -2320
rect 6483 -2429 6564 -2427
rect 3576 -2511 3583 -2455
rect 3639 -2511 3657 -2455
rect 9105 -2477 9181 -2376
rect 9333 -2322 9409 -2312
rect 9333 -2378 9343 -2322
rect 9399 -2378 9409 -2322
rect 10122 -2352 10133 -2296
rect 10189 -2352 11256 -2296
rect 11368 -2352 11424 -2296
rect 10122 -2362 10198 -2352
rect 9333 -2388 9409 -2378
rect 11227 -2381 11396 -2352
rect 3576 -2528 3657 -2511
rect 7556 -2486 9181 -2477
rect 7556 -2538 7573 -2486
rect 7625 -2538 9181 -2486
rect 7556 -2556 9181 -2538
rect 7556 -2557 9171 -2556
rect 3686 -2730 4020 -2710
rect 3686 -2810 3764 -2730
rect 3926 -2810 4020 -2730
rect 3686 -2830 4020 -2810
rect 5649 -2734 5983 -2710
rect 5649 -2814 5724 -2734
rect 5886 -2814 5983 -2734
rect 5649 -2830 5983 -2814
rect 7662 -2730 7996 -2710
rect 7662 -2810 7752 -2730
rect 7914 -2810 7996 -2730
rect 7662 -2830 7996 -2810
<< via2 >>
rect 2838 1329 3000 1409
rect 4573 1333 4735 1413
rect 6674 1332 6836 1412
rect 3768 549 3930 629
rect 5736 553 5898 633
rect 7744 549 7906 629
rect 2828 217 2990 297
rect 4600 213 4762 293
rect 6660 221 6822 301
rect 3772 -571 3934 -491
rect 5744 -567 5906 -487
rect 7752 -567 7914 -487
rect 2852 -903 3014 -823
rect 4584 -911 4746 -831
rect 6664 -903 6826 -823
rect 3768 -1695 3930 -1615
rect 5728 -1687 5890 -1607
rect 7740 -1691 7902 -1611
rect 2836 -2023 2998 -1943
rect 4580 -2027 4742 -1947
rect 6668 -2027 6830 -1947
rect 3764 -2810 3926 -2730
rect 5724 -2814 5886 -2734
rect 7752 -2810 7914 -2730
<< metal3 >>
rect 2770 1409 3104 1721
rect 2770 1329 2838 1409
rect 3000 1329 3104 1409
rect 2770 297 3104 1329
rect 2770 217 2828 297
rect 2990 217 3104 297
rect 2770 -199 3104 217
rect 2770 -279 2855 -199
rect 3017 -279 3104 -199
rect 2770 -823 3104 -279
rect 2770 -903 2852 -823
rect 3014 -903 3104 -823
rect 2770 -1723 3104 -903
rect 2770 -1803 2845 -1723
rect 3007 -1803 3104 -1723
rect 2770 -1943 3104 -1803
rect 2770 -2023 2836 -1943
rect 2998 -2023 3104 -1943
rect 2770 -2976 3104 -2023
rect 3686 629 4020 1721
rect 3686 549 3768 629
rect 3930 549 4020 629
rect 3686 -491 4020 549
rect 3686 -571 3772 -491
rect 3934 -571 4020 -491
rect 3686 -891 4020 -571
rect 3686 -971 3756 -891
rect 3918 -971 4020 -891
rect 3686 -1615 4020 -971
rect 3686 -1695 3768 -1615
rect 3930 -1695 4020 -1615
rect 3686 -2730 4020 -1695
rect 3686 -2810 3764 -2730
rect 3926 -2810 4020 -2730
rect 3686 -2976 4020 -2810
rect 4508 1413 4842 1672
rect 4508 1333 4573 1413
rect 4735 1333 4842 1413
rect 4508 293 4842 1333
rect 4508 213 4600 293
rect 4762 213 4842 293
rect 4508 -218 4842 213
rect 4508 -298 4574 -218
rect 4736 -298 4842 -218
rect 4508 -831 4842 -298
rect 4508 -911 4584 -831
rect 4746 -911 4842 -831
rect 4508 -1723 4842 -911
rect 4508 -1803 4591 -1723
rect 4753 -1803 4842 -1723
rect 4508 -1947 4842 -1803
rect 4508 -2027 4580 -1947
rect 4742 -2027 4842 -1947
rect 4508 -3025 4842 -2027
rect 5649 633 5983 1666
rect 5649 553 5736 633
rect 5898 553 5983 633
rect 5649 -487 5983 553
rect 5649 -567 5744 -487
rect 5906 -567 5983 -487
rect 5649 -891 5983 -567
rect 5649 -971 5728 -891
rect 5890 -971 5983 -891
rect 5649 -1607 5983 -971
rect 5649 -1687 5728 -1607
rect 5890 -1687 5983 -1607
rect 5649 -2734 5983 -1687
rect 5649 -2814 5724 -2734
rect 5886 -2814 5983 -2734
rect 5649 -3031 5983 -2814
rect 6581 1412 6915 1644
rect 6581 1332 6674 1412
rect 6836 1332 6915 1412
rect 6581 301 6915 1332
rect 6581 221 6660 301
rect 6822 221 6915 301
rect 6581 -250 6915 221
rect 6581 -330 6681 -250
rect 6843 -330 6915 -250
rect 6581 -823 6915 -330
rect 6581 -903 6664 -823
rect 6826 -903 6915 -823
rect 6581 -1724 6915 -903
rect 6581 -1804 6670 -1724
rect 6832 -1804 6915 -1724
rect 6581 -1947 6915 -1804
rect 6581 -2027 6668 -1947
rect 6830 -2027 6915 -1947
rect 6581 -3053 6915 -2027
rect 7662 629 7996 1633
rect 7662 549 7744 629
rect 7906 549 7996 629
rect 7662 -487 7996 549
rect 7662 -567 7752 -487
rect 7914 -567 7996 -487
rect 7662 -903 7996 -567
rect 7662 -983 7738 -903
rect 7900 -983 7996 -903
rect 7662 -1611 7996 -983
rect 7662 -1691 7740 -1611
rect 7902 -1691 7996 -1611
rect 7662 -2730 7996 -1691
rect 7662 -2810 7752 -2730
rect 7914 -2810 7996 -2730
rect 7662 -3064 7996 -2810
<< via3 >>
rect 2838 1329 3000 1409
rect 2855 -279 3017 -199
rect 2845 -1803 3007 -1723
rect 3768 549 3930 629
rect 3756 -971 3918 -891
rect 3764 -2810 3926 -2730
rect 4573 1333 4735 1413
rect 4574 -298 4736 -218
rect 4591 -1803 4753 -1723
rect 5736 553 5898 633
rect 5728 -971 5890 -891
rect 5724 -2814 5886 -2734
rect 6674 1332 6836 1412
rect 6681 -330 6843 -250
rect 6670 -1804 6832 -1724
rect 7744 549 7906 629
rect 7738 -983 7900 -903
rect 7752 -2810 7914 -2730
<< metal4 >>
rect 1844 1413 11646 1505
rect 1844 1409 4573 1413
rect 1844 1329 2838 1409
rect 3000 1333 4573 1409
rect 4735 1412 11646 1413
rect 4735 1333 6674 1412
rect 3000 1332 6674 1333
rect 6836 1332 11646 1412
rect 3000 1329 11646 1332
rect 1844 1170 11646 1329
rect 1838 633 11640 709
rect 1838 629 5736 633
rect 1838 549 3768 629
rect 3930 553 5736 629
rect 5898 629 11640 633
rect 5898 553 7744 629
rect 3930 549 7744 553
rect 7906 549 11640 629
rect 1838 374 11640 549
rect 1868 -199 11670 -80
rect 1868 -279 2855 -199
rect 3017 -218 11670 -199
rect 3017 -279 4574 -218
rect 1868 -298 4574 -279
rect 4736 -250 11670 -218
rect 4736 -298 6681 -250
rect 1868 -330 6681 -298
rect 6843 -330 11670 -250
rect 1868 -415 11670 -330
rect 1874 -891 11676 -780
rect 1874 -971 3756 -891
rect 3918 -971 5728 -891
rect 5890 -903 11676 -891
rect 5890 -971 7738 -903
rect 1874 -983 7738 -971
rect 7900 -983 11676 -903
rect 1874 -1115 11676 -983
rect 1904 -1723 11706 -1576
rect 1904 -1803 2845 -1723
rect 3007 -1803 4591 -1723
rect 4753 -1724 11706 -1723
rect 4753 -1803 6670 -1724
rect 1904 -1804 6670 -1803
rect 6832 -1804 11706 -1724
rect 1904 -1911 11706 -1804
rect 1922 -2730 11724 -2557
rect 1922 -2810 3764 -2730
rect 3926 -2734 7752 -2730
rect 3926 -2810 5724 -2734
rect 1922 -2814 5724 -2810
rect 5886 -2810 7752 -2734
rect 7914 -2810 11724 -2730
rect 5886 -2814 11724 -2810
rect 1922 -2892 11724 -2814
use CS_Switch_1x1  CS_Switch_1x1_0
timestamp 1755764817
transform 1 0 9064 0 1 938
box -306 -434 837 214
use CS_Switch_2x2  CS_Switch_2x2_1
timestamp 1755705199
transform 1 0 9106 0 1 -180
box -356 -436 795 224
use CS_Switch_4x2  CS_Switch_4x2_0
timestamp 1755705775
transform 1 0 9054 0 1 -1551
box -304 -185 1117 488
use CS_Switch_8x2  CS_Switch_8x2_0
timestamp 1755706082
transform 1 0 8387 0 1 -3880
box 426 1024 1804 1719
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 7766 0 1 590
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_1
timestamp 1753044640
transform 1 0 6870 0 1 -2770
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_4
timestamp 1753044640
transform 1 0 6870 0 1 -1650
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_5
timestamp 1753044640
transform 1 0 7766 0 1 -2770
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_6
timestamp 1753044640
transform 1 0 6870 0 1 -530
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_7
timestamp 1753044640
transform 1 0 7766 0 1 -1650
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_8
timestamp 1753044640
transform 1 0 6870 0 1 590
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_9
timestamp 1753044640
transform 1 0 7766 0 1 -530
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2662 0 1 -2770
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_1
timestamp 1753044640
transform 1 0 2662 0 1 590
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_2
timestamp 1753044640
transform 1 0 2662 0 1 -530
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_3
timestamp 1753044640
transform 1 0 2662 0 1 -1650
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 6134 0 1 -530
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_1
timestamp 1753044640
transform 1 0 6134 0 1 590
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_2
timestamp 1753044640
transform 1 0 6134 0 1 -2770
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_3
timestamp 1753044640
transform 1 0 6134 0 1 -1650
box -86 -86 758 870
<< labels >>
flabel metal2 3576 832 3657 1132 1 FreeSans 800 0 0 0 D1
port 1 n
flabel metal2 3576 -288 3657 12 1 FreeSans 800 0 0 0 D2
port 2 n
flabel metal2 3576 -1408 3657 -1108 1 FreeSans 800 0 0 0 D3
port 3 n
flabel metal2 3576 -2528 3657 -2228 1 FreeSans 800 0 0 0 D4
port 4 n
flabel metal3 2770 1409 3104 1721 1 FreeSans 3200 0 0 0 VDD
port 9 n
flabel metal3 3686 629 4020 1721 1 FreeSans 3200 0 0 0 VSS
port 10 n
flabel metal1 10248 -2912 10584 1624 1 FreeSans 800 0 0 0 OUTN
port 6 n
flabel metal1 10696 -2912 11032 1624 1 FreeSans 800 0 0 0 OUTP
port 5 n
flabel metal1 11144 -2912 11480 1624 1 FreeSans 800 0 0 0 VBIAS
port 7 n
flabel metal1 2240 -2968 2576 1680 1 FreeSans 800 0 0 0 CLK
port 8 n
<< properties >>
string CS_Switch_2x2_0 x1
string name x1
<< end >>
