magic
tech gf180mcuD
magscale 1 10
timestamp 1754362338
<< pwell >>
rect 687 856 2281 1496
<< nmos >>
rect 896 1232 952 1276
rect 1124 1233 1180 1277
rect 1489 1232 1545 1276
rect 1637 1208 1997 1296
<< ndiff >>
rect 770 1276 850 1293
rect 998 1277 1078 1294
rect 1226 1277 1306 1294
rect 998 1276 1124 1277
rect 770 1275 896 1276
rect 770 1228 787 1275
rect 833 1232 896 1275
rect 952 1232 1015 1276
rect 833 1228 850 1232
rect 770 1211 850 1228
rect 998 1229 1015 1232
rect 1061 1233 1124 1276
rect 1180 1276 1306 1277
rect 1180 1233 1243 1276
rect 1061 1229 1078 1233
rect 998 1212 1078 1229
rect 1226 1229 1243 1233
rect 1289 1229 1306 1276
rect 1226 1212 1306 1229
rect 1363 1276 1443 1294
rect 1591 1276 1637 1296
rect 1363 1229 1380 1276
rect 1426 1232 1489 1276
rect 1545 1232 1637 1276
rect 1426 1229 1443 1232
rect 1363 1212 1443 1229
rect 1591 1208 1637 1232
rect 1997 1293 2043 1296
rect 1997 1275 2123 1293
rect 1997 1228 2060 1275
rect 2106 1228 2123 1275
rect 1997 1211 2123 1228
rect 1997 1208 2043 1211
<< ndiffc >>
rect 787 1228 833 1275
rect 1015 1229 1061 1276
rect 1243 1229 1289 1276
rect 1380 1229 1426 1276
rect 2060 1228 2106 1275
<< polysilicon >>
rect 885 1386 965 1404
rect 885 1340 901 1386
rect 947 1340 965 1386
rect 885 1322 965 1340
rect 1113 1387 1193 1405
rect 1113 1341 1129 1387
rect 1175 1341 1193 1387
rect 1113 1323 1193 1341
rect 1488 1378 1997 1400
rect 1488 1332 1765 1378
rect 1885 1332 1997 1378
rect 896 1276 952 1322
rect 1124 1277 1180 1323
rect 1488 1316 1997 1332
rect 896 1186 952 1232
rect 1124 1187 1180 1233
rect 1489 1276 1545 1316
rect 1637 1296 1997 1316
rect 1489 1186 1545 1232
rect 1637 1163 1997 1208
<< polycontact >>
rect 901 1340 947 1386
rect 1129 1341 1175 1387
rect 1765 1332 1885 1378
<< metal1 >>
rect 781 1290 837 1449
rect 896 1386 952 1449
rect 896 1340 901 1386
rect 947 1340 952 1386
rect 896 1329 952 1340
rect 1124 1387 1180 1450
rect 1124 1341 1129 1387
rect 1175 1341 1180 1387
rect 1124 1330 1180 1341
rect 1237 1291 1293 1448
rect 1690 1378 1953 1391
rect 1690 1332 1765 1378
rect 1885 1332 1953 1378
rect 1690 1320 1953 1332
rect 772 1275 848 1290
rect 772 1228 787 1275
rect 833 1228 848 1275
rect 772 1213 848 1228
rect 1000 1276 1076 1291
rect 1000 1229 1015 1276
rect 1061 1229 1076 1276
rect 1000 1214 1076 1229
rect 1228 1276 1304 1291
rect 1228 1229 1243 1276
rect 1289 1229 1304 1276
rect 1228 1214 1304 1229
rect 1365 1276 1441 1291
rect 1365 1229 1380 1276
rect 1426 1229 1441 1276
rect 1365 1214 1441 1229
rect 2045 1275 2121 1290
rect 2045 1228 2060 1275
rect 2106 1228 2121 1275
rect 1008 1162 1064 1214
rect 1376 1162 1432 1214
rect 2045 1213 2121 1228
rect 1007 1106 1432 1162
rect 2056 1043 2112 1213
rect 1886 1042 2219 1043
rect 772 951 2219 1042
<< labels >>
flabel metal1 900 1334 948 1438 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 1128 1336 1176 1440 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 784 1222 836 1420 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 1239 1223 1291 1421 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 1724 1327 1934 1389 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 2059 1001 2111 1286 1 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional
flabel pwell 783 958 1044 1030 1 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
<< end >>
