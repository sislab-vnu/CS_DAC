magic
tech gf180mcuD
magscale 1 10
timestamp 1754652878
<< pwell >>
rect 4495 -2762 4890 -2693
rect 4904 -2762 4973 -2367
rect 3723 -3319 3969 -3111
<< metal1 >>
rect 3414 -348 3656 783
rect 3764 -301 3793 -237
rect 3901 -301 5062 -237
rect 4998 -302 5062 -301
rect 3414 -412 4651 -348
rect 3414 -413 3657 -412
rect 3414 -1208 3656 -413
rect 4589 -682 4651 -412
rect 4998 -609 5063 -302
rect 9660 -513 9736 -512
rect 4972 -674 5063 -609
rect 5983 -602 6312 -519
rect 9441 -589 9736 -513
rect 5200 -1001 5447 -883
rect 3414 -1273 3657 -1208
rect 3789 -1224 3801 -1160
rect 3910 -1224 5037 -1160
rect 3414 -1337 4626 -1273
rect 3414 -2225 3657 -1337
rect 4563 -1599 4626 -1337
rect 4975 -1362 5037 -1224
rect 4974 -1599 5037 -1362
rect 9660 -1469 9736 -589
rect 5989 -1558 6309 -1475
rect 9457 -1546 9736 -1469
rect 5237 -1959 5446 -1839
rect 5237 -1960 5319 -1959
rect 3777 -2117 4780 -2116
rect 3777 -2179 3792 -2117
rect 3902 -2179 4780 -2117
rect 4719 -2212 4780 -2179
rect 3414 -2289 4374 -2225
rect 3414 -3449 3657 -2289
rect 4311 -2554 4374 -2289
rect 4719 -2554 4782 -2287
rect 9660 -2432 9736 -1546
rect 5986 -2521 6326 -2438
rect 9456 -2508 9736 -2432
rect 5210 -2922 5498 -2802
rect 3783 -3309 3802 -3247
rect 3898 -3248 4743 -3247
rect 3898 -3308 4913 -3248
rect 3898 -3309 4269 -3308
rect 4741 -3309 4913 -3308
rect 3414 -3450 4008 -3449
rect 3414 -3514 4541 -3450
rect 3414 -3515 4008 -3514
rect 3414 -3530 3657 -3515
rect 4852 -3517 4913 -3309
rect 9660 -3404 9736 -2508
rect 5989 -3493 6327 -3410
rect 9456 -3480 9736 -3404
rect 9660 -3570 9736 -3480
rect 5232 -3894 5451 -3774
<< via1 >>
rect 3793 -301 3901 -237
rect 4407 -548 4463 -496
rect 4711 -547 4765 -494
rect 4878 -548 4936 -494
rect 6341 -460 6481 -374
rect 5581 -634 5641 -547
rect 3801 -1224 3910 -1160
rect 4384 -1464 4437 -1412
rect 4686 -1466 4741 -1413
rect 4863 -1467 4917 -1413
rect 6351 -1406 6474 -1340
rect 5581 -1590 5641 -1505
rect 3792 -2179 3902 -2117
rect 4128 -2420 4181 -2368
rect 4429 -2421 4484 -2367
rect 4606 -2421 4661 -2367
rect 4911 -2420 4965 -2367
rect 6357 -2371 6473 -2302
rect 5582 -2554 5642 -2470
rect 3802 -3309 3898 -3247
rect 4594 -3422 4651 -3369
rect 4736 -3423 4793 -3370
rect 6361 -3341 6475 -3281
rect 5582 -3524 5642 -3437
rect 4383 -3625 4438 -3572
rect 4950 -3624 5003 -3571
<< metal2 >>
rect 3717 287 3968 781
rect 3717 -237 3969 287
rect 3717 -301 3793 -237
rect 3901 -301 3969 -237
rect 3717 -606 3969 -301
rect 4037 -484 4280 781
rect 4701 -355 5457 -354
rect 6305 -355 6521 -348
rect 4701 -374 6521 -355
rect 4701 -423 6341 -374
rect 4701 -481 4780 -423
rect 5001 -424 6341 -423
rect 6305 -460 6341 -424
rect 6481 -460 6521 -374
rect 6305 -477 6521 -460
rect 4395 -484 4475 -481
rect 4037 -496 4475 -484
rect 4037 -548 4407 -496
rect 4463 -548 4475 -496
rect 4037 -559 4475 -548
rect 3717 -617 3968 -606
rect 3720 -737 3968 -617
rect 3720 -1160 3969 -737
rect 3720 -1224 3801 -1160
rect 3910 -1224 3969 -1160
rect 3720 -2117 3969 -1224
rect 3720 -2162 3792 -2117
rect 3723 -2179 3792 -2162
rect 3902 -2179 3969 -2117
rect 3723 -2218 3969 -2179
rect 3722 -3247 3969 -2218
rect 3722 -3309 3802 -3247
rect 3898 -3309 3969 -3247
rect 3722 -3319 3969 -3309
rect 4037 -1402 4280 -559
rect 4395 -561 4475 -559
rect 4699 -494 4780 -481
rect 4699 -547 4711 -494
rect 4765 -508 4780 -494
rect 4867 -490 4947 -481
rect 4867 -494 5662 -490
rect 4765 -547 4779 -508
rect 4699 -561 4779 -547
rect 4867 -548 4878 -494
rect 4936 -547 5662 -494
rect 4936 -548 5581 -547
rect 4867 -559 5581 -548
rect 4867 -561 4947 -559
rect 5551 -634 5581 -559
rect 5641 -559 5662 -547
rect 5641 -634 5661 -559
rect 5551 -648 5661 -634
rect 4675 -1340 6524 -1271
rect 4675 -1341 6351 -1340
rect 4675 -1399 4751 -1341
rect 4370 -1402 4450 -1399
rect 4037 -1412 4450 -1402
rect 4037 -1464 4384 -1412
rect 4437 -1464 4450 -1412
rect 4037 -1477 4450 -1464
rect 4037 -2368 4280 -1477
rect 4370 -1479 4450 -1477
rect 4674 -1413 4754 -1399
rect 4674 -1466 4686 -1413
rect 4741 -1466 4754 -1413
rect 4674 -1479 4754 -1466
rect 4850 -1409 4930 -1399
rect 6307 -1406 6351 -1341
rect 6474 -1341 6524 -1340
rect 6474 -1406 6523 -1341
rect 4850 -1413 5663 -1409
rect 4850 -1467 4863 -1413
rect 4917 -1467 5663 -1413
rect 6307 -1433 6523 -1406
rect 4850 -1479 5663 -1467
rect 5555 -1505 5663 -1479
rect 5555 -1590 5581 -1505
rect 5641 -1590 5663 -1505
rect 5555 -1604 5663 -1590
rect 4419 -2159 6523 -2089
rect 4419 -2354 4486 -2159
rect 4596 -2290 5640 -2220
rect 4596 -2354 4672 -2290
rect 4037 -2420 4128 -2368
rect 4181 -2420 4280 -2368
rect 4037 -2693 4280 -2420
rect 4418 -2367 4498 -2354
rect 4418 -2421 4429 -2367
rect 4484 -2421 4498 -2367
rect 4418 -2434 4498 -2421
rect 4594 -2367 4674 -2354
rect 4594 -2421 4606 -2367
rect 4661 -2421 4674 -2367
rect 4594 -2434 4674 -2421
rect 4898 -2367 4978 -2354
rect 4898 -2420 4911 -2367
rect 4965 -2420 4978 -2367
rect 4898 -2434 4978 -2420
rect 4904 -2693 4973 -2434
rect 5555 -2449 5640 -2290
rect 6308 -2267 6523 -2159
rect 6308 -2302 6524 -2267
rect 6308 -2371 6357 -2302
rect 6473 -2371 6524 -2302
rect 6308 -2396 6524 -2371
rect 5555 -2470 5669 -2449
rect 5555 -2554 5582 -2470
rect 5642 -2554 5669 -2470
rect 5555 -2567 5669 -2554
rect 5555 -2568 5666 -2567
rect 4037 -2762 4973 -2693
rect 3722 -3412 3968 -3319
rect 4037 -3563 4280 -2762
rect 4585 -3281 6524 -3219
rect 4585 -3289 6361 -3281
rect 4585 -3356 4656 -3289
rect 6308 -3341 6361 -3289
rect 6475 -3341 6524 -3281
rect 4584 -3369 4664 -3356
rect 4584 -3422 4594 -3369
rect 4651 -3422 4664 -3369
rect 4584 -3436 4664 -3422
rect 4724 -3365 4804 -3356
rect 4724 -3370 5665 -3365
rect 6308 -3368 6524 -3341
rect 4724 -3423 4736 -3370
rect 4793 -3423 5665 -3370
rect 4724 -3435 5665 -3423
rect 4724 -3436 4804 -3435
rect 5558 -3437 5664 -3435
rect 5558 -3524 5582 -3437
rect 5642 -3524 5664 -3437
rect 5558 -3539 5664 -3524
rect 4372 -3563 4452 -3558
rect 4037 -3564 4452 -3563
rect 4936 -3564 5016 -3558
rect 4037 -3571 5016 -3564
rect 4037 -3572 4950 -3571
rect 4037 -3625 4383 -3572
rect 4438 -3624 4950 -3572
rect 5003 -3624 5016 -3571
rect 4438 -3625 5016 -3624
rect 4037 -3634 5016 -3625
rect 4037 -3636 4452 -3634
rect 4037 -3658 4280 -3636
rect 4372 -3638 4452 -3636
rect 4936 -3638 5016 -3634
use CS_Switch_1x1  CS_Switch_1x1_0
timestamp 1754553491
transform -1 0 4935 0 1 -627
box -382 -434 929 214
use CS_Switch_2x2  CS_Switch_2x2_0
timestamp 1754556308
transform -1 0 4894 0 1 -1563
box -438 -436 877 224
use CS_Switch_4x2  CS_Switch_4x2_0
timestamp 1754559251
transform 1 0 4140 0 1 -2778
box -376 -185 1183 488
use CS_Switch_8x2  CS_Switch_8x2_0
timestamp 1754627642
transform 1 0 3556 0 1 -5460
box 518 1526 1757 2149
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform -1 0 9590 0 1 -2862
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_1
timestamp 1753044640
transform -1 0 9587 0 1 -943
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_2
timestamp 1753044640
transform -1 0 9589 0 1 -1899
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_3
timestamp 1753044640
transform -1 0 9590 0 1 -3834
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform -1 0 6118 0 1 -2862
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_1
timestamp 1753044640
transform -1 0 6117 0 1 -943
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_2
timestamp 1753044640
transform -1 0 6117 0 1 -1899
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_3
timestamp 1753044640
transform -1 0 6118 0 1 -3834
box -86 -86 758 870
<< labels >>
flabel space 8592 -701 8673 -401 1 FreeSans 400 0 0 0 D1
port 1 n
flabel space 8594 -1657 8675 -1357 1 FreeSans 400 0 0 0 D2
port 2 n
flabel space 8595 -2620 8676 -2320 1 FreeSans 400 0 0 0 D3
port 3 n
flabel space 8595 -3592 8676 -3292 1 FreeSans 400 0 0 0 D4
port 4 n
flabel metal1 9660 -3570 9736 -512 1 FreeSans 400 0 0 0 CLK
port 5 n
flabel metal1 3414 -3530 3656 783 1 FreeSans 400 0 0 0 OUTP
port 6 n
flabel metal2 3720 -2117 3969 -1224 1 FreeSans 400 0 0 0 OUTN
port 7 n
flabel metal2 4037 -2368 4280 781 1 FreeSans 400 0 0 0 VBIAS
port 8 n
<< end >>
