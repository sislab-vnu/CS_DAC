* NGSPICE file created from CS_Switch_1x.ext - technology: gf180mcuD

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT layouted_cell__CS_Switch_1x INP INN OUTP OUTN VBIAS VSS VPW
X0 a_668_n40# VSS a_440_n224# VPW nfet_03v3 ad=50.6f pd=0.9u as=0.1452p ps=1.465u w=0.22u l=0.28u
X1 a_668_n224# VSS a_440_n224# VPW nfet_03v3 ad=50.6f pd=0.9u as=0.1452p ps=1.465u w=0.22u l=0.28u
X2 a_440_n224# VBIAS a_56_n40# VPW nfet_03v3 ad=0.1452p pd=1.465u as=0.1516p ps=1.64u w=0.22u l=0.28u
X3 VSS VSS a_n228_n224# VPW nfet_03v3 ad=94.5f pd=0.99u as=50.6f ps=0.9u w=0.22u l=0.28u
X4 OUTN INN a_56_n40# VPW nfet_03v3 ad=0.182p pd=1.8u as=86.8f ps=0.92u w=0.22u l=0.28u
X5 a_440_n224# VBIAS VSS VPW nfet_03v3 ad=0.1452p pd=1.465u as=94.5f ps=0.99u w=0.22u l=2.2u
X6 a_56_n40# INP OUTP VPW nfet_03v3 ad=86.8f pd=0.92u as=0.1053p ps=1.03u w=0.22u l=0.28u
X7 OUTP VSS a_n228_n40# VPW nfet_03v3 ad=0.1053p pd=1.03u as=50.6f ps=0.9u w=0.22u l=0.28u
C0 a_440_n224# VSS 0.006325f
C1 VPW INP 0.105738f
C2 a_n228_n224# VSS 3.61e-19
C3 a_440_n224# VBIAS 0.001013f
C4 INN VBIAS 0.041164f
C5 OUTN INP 7.62e-20
C6 VPW VSS 0.275976f
C7 OUTN VSS 4.68e-20
C8 VSS a_n228_n40# 2.43e-19
C9 VPW VBIAS 0.410847f
C10 VSS a_668_n40# 5.59e-19
C11 OUTN VBIAS 0.001717f
C12 VSS a_668_n224# 8.29e-19
C13 VSS INP 0.021464f
C14 INP VBIAS 0.019271f
C15 OUTP a_56_n40# 0.029701f
C16 VSS VBIAS 0.11846f
C17 OUTP INN 7.62e-20
C18 a_440_n224# a_56_n40# 0.00171f
C19 INN a_56_n40# 0.029406f
C20 OUTN OUTP 6.32e-19
C21 a_n228_n40# OUTP 7.7e-19
C22 OUTN a_56_n40# 0.164087f
C23 VPW INN 0.108806f
C24 INP OUTP 0.003858f
C25 OUTN INN 0.003858f
C26 INP a_56_n40# 0.003069f
C27 VSS OUTP 0.02973f
C28 VSS a_56_n40# 0.150521f
C29 a_56_n40# VBIAS 0.047893f
C30 INP INN 0.060872f
C31 OUTN VSUBS 0.018808f
C32 OUTP VSUBS 0.030912f
C33 VSS VSUBS 0.66916f
C34 VBIAS VSUBS 0.414038f
C35 INN VSUBS 0.069304f
C36 INP VSUBS 0.085275f
C37 a_56_n40# VSUBS 0.105866f
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT layouted_cell__CS_Switch_2x INP INN OUTP OUTN VBIAS VSS VPW
X0 a_n226_n248# VSS a_n328_n248# VPW nfet_03v3 ad=0.1012p pd=1.34u as=0.1012p ps=1.34u w=0.44u l=0.28u
X1 a_n226_n20# VSS a_n366_n20# VPW nfet_03v3 ad=50.6f pd=0.9u as=92.4f ps=1.28u w=0.22u l=0.28u
X2 a_336_n248# VBIAS a_32_n20# VPW nfet_03v3 ad=0.2695p pd=2.66u as=0.1516p ps=1.64u w=0.22u l=0.28u
X3 OUTN INN a_32_n20# VPW nfet_03v3 ad=0.182p pd=1.8u as=0.102p ps=1u w=0.22u l=0.28u
X4 a_734_n20# VSS a_632_n20# VPW nfet_03v3 ad=92.4f pd=1.28u as=50.6f ps=0.9u w=0.22u l=0.28u
X5 a_32_n20# INP OUTP VPW nfet_03v3 ad=0.102p pd=1u as=0.182p ps=1.8u w=0.22u l=0.28u
X6 a_336_n248# VBIAS VSS VPW nfet_03v3 ad=0.2695p pd=2.66u as=0.1932p ps=1.8u w=0.44u l=1.8u
X7 a_734_n248# VSS a_632_n248# VPW nfet_03v3 ad=0.1012p pd=1.34u as=0.1012p ps=1.34u w=0.44u l=0.28u
C0 OUTP VSS 0.026879f
C1 a_n366_n20# VSS 7.12e-19
C2 a_734_n20# VSS 7.12e-19
C3 VBIAS INN 0.041085f
C4 OUTP INN 7.31e-20
C5 VSS a_336_n248# 0.009017f
C6 OUTN INP 7.31e-20
C7 a_32_n20# VBIAS 0.049088f
C8 VSS a_n226_n248# 0.003027f
C9 a_32_n20# OUTP 0.028781f
C10 VSS OUTN 3.28e-20
C11 a_n226_n20# VSS 4.96e-19
C12 VSS INP 0.016517f
C13 a_n366_n20# OUTP 0.001129f
C14 OUTN INN 0.003859f
C15 a_32_n20# a_336_n248# 0.004061f
C16 INN INP 0.055413f
C17 VBIAS a_336_n248# 0.001019f
C18 a_n328_n248# VSS 0.002749f
C19 a_32_n20# OUTN 0.163167f
C20 VSS a_632_n20# 4.96e-19
C21 a_32_n20# INP 0.003036f
C22 VSS a_632_n248# 0.001897f
C23 VBIAS OUTN 0.001721f
C24 OUTP OUTN 6.13e-19
C25 a_734_n248# VSS 0.00184f
C26 VBIAS INP 0.019794f
C27 a_n226_n20# OUTP 8.03e-19
C28 OUTP INP 0.003859f
C29 a_32_n20# VSS 0.10817f
C30 VBIAS VSS 0.109396f
C31 a_32_n20# INN 0.029571f
C32 OUTN VPW 0.018761f
C33 OUTP VPW 0.030882f
C34 VSS VPW 1.06828f
C35 VBIAS VPW 0.790242f
C36 INN VPW 0.178433f
C37 INP VPW 0.194214f
C38 a_32_n20# VPW 0.108528f
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT layouted_cell__CS_Switch_4x INP INN OUTP OUTN VBIAS VSS VPW
X0 a_1050_0# VSS a_948_0# VPW nfet_03v3 ad=0.1035p pd=1.36u as=0.1035p ps=1.36u w=0.45u l=0.28u
X1 a_42_240# INP OUTP VPW nfet_03v3 ad=0.102p pd=1u as=0.182p ps=1.8u w=0.22u l=0.28u
X2 a_812_0# VBIAS a_42_240# VPW nfet_03v3 ad=0.21255p pd=1.92u as=0.1516p ps=1.64u w=0.22u l=0.28u
X3 VSS VBIAS a_n80_0# VPW nfet_03v3 ad=0.2128p pd=1.78u as=0.21255p ps=1.92u w=0.45u l=1.8u
X4 a_42_240# VBIAS a_n80_0# VPW nfet_03v3 ad=0.1516p pd=1.64u as=0.21255p ps=1.92u w=0.22u l=0.28u
X5 OUTN INN a_42_240# VPW nfet_03v3 ad=0.182p pd=1.8u as=0.102p ps=1u w=0.22u l=0.28u
X6 a_n182_0# VSS a_n284_0# VPW nfet_03v3 ad=0.1035p pd=1.36u as=0.1035p ps=1.36u w=0.45u l=0.28u
X7 a_1050_240# VSS a_948_240# VPW nfet_03v3 ad=92.4f pd=1.28u as=50.6f ps=0.9u w=0.22u l=0.28u
X8 a_812_0# VBIAS VSS VPW nfet_03v3 ad=0.21255p pd=1.92u as=0.2128p ps=1.78u w=0.45u l=1.8u
X9 a_n182_240# VSS a_n322_240# VPW nfet_03v3 ad=50.6f pd=0.9u as=92.4f ps=1.28u w=0.22u l=0.28u
C0 a_812_0# VBIAS 6.69e-19
C1 a_812_0# VSS 0.005768f
C2 OUTP INP 0.003859f
C3 OUTN INP 3.66e-20
C4 VSS a_n182_0# 0.001662f
C5 a_42_240# OUTP 0.145304f
C6 a_42_240# OUTN 0.145304f
C7 VBIAS INP 0.038981f
C8 a_42_240# VBIAS 0.096115f
C9 a_948_0# VSS 0.001662f
C10 a_1050_240# VSS 3.37e-19
C11 a_42_240# VSS 0.205235f
C12 a_n322_240# VSS 3.58e-19
C13 VSS a_n182_240# 4.85e-19
C14 a_42_240# a_n80_0# 0.00195f
C15 OUTP OUTN 3.07e-19
C16 OUTP VBIAS 0.001662f
C17 VBIAS OUTN 0.001662f
C18 OUTP VSS 3.26e-20
C19 OUTN VSS 3.26e-20
C20 VBIAS VSS 0.170383f
C21 VSS a_n284_0# 0.001229f
C22 VBIAS a_n80_0# 6.69e-19
C23 a_n80_0# VSS 0.005768f
C24 INN INP 0.055413f
C25 a_42_240# INN 0.028229f
C26 VSS a_948_240# 4.85e-19
C27 a_42_240# a_812_0# 0.00195f
C28 a_42_240# INP 0.028229f
C29 OUTP INN 3.66e-20
C30 OUTN INN 0.003859f
C31 VBIAS INN 0.038981f
C32 a_1050_0# VSS 0.001156f
C33 OUTN VPW 0.019015f
C34 OUTP VPW 0.019015f
C35 VSS VPW 1.05553f
C36 INN VPW 0.179143f
C37 INP VPW 0.179143f
C38 VBIAS VPW 1.4513f
C39 a_42_240# VPW 0.176002f
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT layouted_cell__CS_Switch_8x INP INN OUTP OUTN VBIAS VSS VPW
X0 a_784_1400# INP OUTP VPW nfet_03v3 ad=0.1306p pd=1.26u as=0.1328p ps=1.28u w=0.22u l=0.28u
X1 OUTP VSS a_450_1400# VPW nfet_03v3 ad=0.1328p pd=1.28u as=50.6f ps=0.9u w=0.22u l=0.28u
X2 OUTN INN a_784_1400# VPW nfet_03v3 ad=0.2106p pd=2.06u as=0.1306p ps=1.26u w=0.22u l=0.28u
X3 VSS VBIAS a_1348_1366# VPW nfet_03v3 ad=0.2026p pd=1.6u as=0.1357p ps=1.08u w=0.62u l=0.3u
X4 a_1348_1366# VBIAS a_784_1400# VPW nfet_03v3 ad=0.1357p pd=1.08u as=0.2248p ps=2.06u w=0.56u l=0.28u
X5 a_1712_1360# VSS VSS VPW nfet_03v3 ad=0.1426p pd=1.7u as=0.2026p ps=1.6u w=0.62u l=0.3u
C0 INN OUTN 0.003587f
C1 INP INN 0.034564f
C2 a_784_1400# INN 0.032405f
C3 INP VSS 0.022774f
C4 a_784_1400# VSS 0.445348f
C5 INN VSS 0.001406f
C6 VBIAS a_1348_1366# 0.004224f
C7 VSS a_450_1400# 5.26e-19
C8 a_784_1400# a_1348_1366# 0.003294f
C9 VSS a_1712_1360# 0.003417f
C10 VBIAS INP 1.33e-20
C11 VBIAS a_784_1400# 0.010206f
C12 a_1348_1366# VSS 0.006681f
C13 INP OUTP 0.003587f
C14 a_784_1400# OUTP 0.023319f
C15 VBIAS INN 0.013345f
C16 VBIAS VSS 0.055613f
C17 VSS OUTP 0.026376f
C18 a_784_1400# OUTN 0.154807f
C19 OUTP a_450_1400# 7.35e-19
C20 INP a_784_1400# 0.004996f
C21 OUTN VPW 0.018986f
C22 OUTP VPW 0.031901f
C23 VSS VPW 0.978803f
C24 VBIAS VPW 0.3659f
C25 INN VPW 0.19646f
C26 INP VPW 0.203821f
C27 a_784_1400# VPW 0.115832f
.ENDS


******* EOF

* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT layouted_cell__CS_Switch_16x INP INN OUTP OUTN VBIAS VSS VPW
X0 a_186_832# VBIAS a_64_826# VPW nfet_03v3 ad=0.1763p pd=1.32u as=99.299995f ps=0.95u w=0.56u l=0.28u
X1 a_64_826# VBIAS VSS VPW nfet_03v3 ad=99.299995f pd=0.95u as=0.1958p ps=1.6u w=0.62u l=0.3u
X2 a_334_832# VBIAS a_186_832# VPW nfet_03v3 ad=99.299995f pd=0.95u as=0.1763p ps=1.32u w=0.56u l=0.28u
X3 a_668_826# VSS VSS VPW nfet_03v3 ad=0.1426p pd=1.7u as=0.1958p ps=1.6u w=0.62u l=0.3u
X4 OUTN INN a_186_832# VPW nfet_03v3 ad=0.405p pd=1.95u as=0.23505p ps=1.76u w=0.6u l=0.3u
X5 VSS VBIAS a_334_832# VPW nfet_03v3 ad=0.1958p pd=1.6u as=99.299995f ps=0.95u w=0.62u l=0.3u
X6 a_668_1100# VSS OUTN VPW nfet_03v3 ad=0.138p pd=1.66u as=0.405p ps=1.95u w=0.6u l=0.3u
X7 VSS VSS a_n250_826# VPW nfet_03v3 ad=0.1958p pd=1.6u as=0.1426p ps=1.7u w=0.62u l=0.3u
X8 a_186_832# INP OUTP VPW nfet_03v3 ad=0.23505p pd=1.76u as=0.405p ps=1.95u w=0.6u l=0.3u
X9 OUTP VSS a_n250_1100# VPW nfet_03v3 ad=0.405p pd=1.95u as=0.138p ps=1.66u w=0.6u l=0.3u
C0 a_186_832# INP 5.25e-19
C1 INN VSS 0.013256f
C2 OUTP VSS 0.013391f
C3 a_186_832# OUTN 0.002131f
C4 OUTP INN 0.001145f
C5 OUTN a_668_1100# 0.001132f
C6 OUTN INP 0.001145f
C7 a_668_826# VSS 0.003029f
C8 a_186_832# VBIAS 0.002221f
C9 a_64_826# INP 2.43e-19
C10 VBIAS INP 0.020299f
C11 OUTN VBIAS 0.029999f
C12 a_186_832# VSS 0.010381f
C13 a_668_1100# VSS 0.001094f
C14 INN a_186_832# 5.25e-19
C15 OUTP a_186_832# 0.002131f
C16 VSS INP 0.013256f
C17 INN INP 0.073624f
C18 OUTP INP 0.002809f
C19 OUTN VSS 0.013391f
C20 a_334_832# VSS 0.004835f
C21 INN OUTN 0.002809f
C22 OUTP OUTN 0.010625f
C23 a_n250_826# VSS 0.003029f
C24 a_334_832# INN 2.43e-19
C25 a_n250_1100# VSS 0.001094f
C26 OUTP a_n250_1100# 0.001132f
C27 a_64_826# VSS 0.004835f
C28 VBIAS VSS 0.140688f
C29 INN VBIAS 0.020299f
C30 OUTP VBIAS 0.029999f
C31 VBIAS VPW 0.630953f
C32 OUTN VPW 0.026697f
C33 OUTP VPW 0.026697f
C34 VSS VPW 1.06007f
C35 INN VPW 0.185395f
C36 INP VPW 0.185395f
.ENDS


******* EOF
