magic
tech gf180mcuD
magscale 1 10
timestamp 1758622440
<< polysilicon >>
rect 157080 112560 157304 128856
rect 157528 112560 157752 128856
rect 157976 112560 158200 128856
rect 158424 112560 158648 128856
rect 158872 112560 159096 128856
rect 159320 112560 159544 128856
rect 159712 112560 159936 128856
rect 160102 128517 176398 128741
rect 185362 128519 200258 128741
rect 160106 128075 176402 128299
rect 185361 128069 200257 128291
rect 160102 127623 176398 127847
rect 185346 127569 200242 127791
rect 160104 127178 176400 127402
rect 185361 127106 200257 127328
rect 160104 126728 176400 126952
rect 185372 126553 200268 126775
rect 160103 126280 176399 126504
rect 185367 126121 200263 126343
rect 160104 125832 176400 126056
rect 185361 125663 200257 125885
rect 160104 125384 176400 125608
rect 185356 125216 200252 125438
rect 160103 124935 176399 125159
rect 185356 124758 200252 124980
rect 160105 124488 176401 124712
rect 156464 94304 156688 105616
rect 156912 94316 157136 105615
rect 157304 94304 157528 105616
rect 157696 94304 157920 105616
rect 158088 94304 158312 105616
rect 158480 94304 158704 105616
rect 158872 94304 159096 105616
rect 159264 94304 159488 105616
rect 159656 94304 159880 105616
rect 160048 94304 160272 98056
rect 160496 94304 160720 98056
<< metal1 >>
rect 156464 112448 156632 132552
rect 159656 112446 159824 132552
rect 176904 124768 177072 132552
rect 180600 127792 180768 132552
rect 176904 124600 177403 124768
rect 188664 123928 188832 132552
rect 212352 128408 212688 132552
rect 212800 128408 213136 132552
rect 213248 128408 213584 132552
rect 160831 123592 204681 123928
rect 212352 123814 212688 123928
rect 212800 123812 213136 123926
rect 213248 123810 213584 123924
<< metal2 >>
rect 154952 94248 156352 129236
rect 156800 112448 156968 132552
rect 157046 128968 184571 130368
rect 157080 112560 157304 128856
rect 157528 112560 157752 128856
rect 157976 112560 158200 128856
rect 158424 112560 158648 128856
rect 158872 112560 159096 128856
rect 159320 112560 159544 128856
rect 159712 112560 159936 128856
rect 160102 128517 176398 128741
rect 160106 128075 176402 128299
rect 160102 127623 176398 127847
rect 184800 127624 184968 132552
rect 185220 128968 200466 130368
rect 185362 128519 200258 128741
rect 185361 128069 200257 128291
rect 184056 127456 184968 127624
rect 185346 127569 200242 127791
rect 160104 127178 176400 127402
rect 185361 127106 200257 127328
rect 160104 126728 176400 126952
rect 160103 126280 176399 126504
rect 160104 125832 176400 126056
rect 160104 125384 176400 125608
rect 160103 124935 176399 125159
rect 160105 124488 176401 124712
rect 177744 124432 177912 125502
rect 161560 124264 177912 124432
rect 161560 123730 161728 124264
rect 178752 124152 178864 126280
rect 167888 123984 178864 124152
rect 167888 123740 168056 123984
rect 179591 123872 179760 125616
rect 174216 123704 179760 123872
rect 180544 123743 180668 126625
rect 181384 123872 181552 125504
rect 182280 124152 182448 126619
rect 185372 126553 200268 126775
rect 185367 126121 200263 126343
rect 183176 124432 183344 125664
rect 185361 125663 200257 125885
rect 185356 125216 200252 125438
rect 185356 124758 200252 124980
rect 200536 124488 200704 132552
rect 200768 128968 202134 130368
rect 202328 125608 202496 132552
rect 202688 128966 203581 130367
rect 203728 126728 203896 132552
rect 204006 128971 205525 130365
rect 205632 127624 205800 132552
rect 205999 128968 215320 130368
rect 203728 126504 205760 126728
rect 202328 125440 205747 125608
rect 183176 124264 199696 124432
rect 200536 124320 205713 124488
rect 182280 123984 193368 124152
rect 181384 123704 187040 123872
rect 193200 123558 193368 123984
rect 199528 123629 199696 124264
rect 160048 119672 161354 119896
rect 160048 111720 160216 119672
rect 158806 111552 160216 111720
rect 160328 116088 161447 116312
rect 160328 110824 160496 116088
rect 157805 110656 160496 110824
rect 160608 112504 161353 112728
rect 160608 109928 160776 112504
rect 158920 109760 160776 109928
rect 157799 108920 161448 109052
rect 158808 107968 160776 108136
rect 158144 107128 160496 107240
rect 158922 106176 160216 106288
rect 156464 94304 156688 105616
rect 156912 94316 157136 105615
rect 157304 94304 157528 105616
rect 157696 94304 157920 105616
rect 158088 94304 158312 105616
rect 158480 94304 158704 105616
rect 158872 94304 159096 105616
rect 159264 94304 159488 105616
rect 159656 94304 159880 105616
rect 160048 98392 160216 106176
rect 160328 101976 160496 107128
rect 160608 105560 160776 107968
rect 160608 105336 161252 105560
rect 160328 101752 161336 101976
rect 160048 98168 161496 98392
rect 160048 94304 160272 98056
rect 160496 94304 160720 98056
rect 213920 94248 215320 128968
rect 154952 93960 215320 94248
rect 154952 93851 214245 93960
rect 156044 92848 214245 93851
<< metal3 >>
rect 152600 132053 154000 132384
rect 152600 131298 152901 132053
rect 153682 131298 154000 132053
rect 152600 121650 154000 131298
rect 215880 132018 217280 132384
rect 215880 131263 216237 132018
rect 217018 131263 217280 132018
rect 154952 130019 215320 130368
rect 154952 129991 214286 130019
rect 154952 129236 155290 129991
rect 156071 129264 214286 129991
rect 215067 129264 215320 130019
rect 156071 129236 215320 129264
rect 154952 128968 215320 129236
rect 162310 123868 162654 128968
rect 163602 123868 163946 128968
rect 165059 123869 165403 128968
rect 168638 123868 168982 128968
rect 169930 123868 170274 128968
rect 171387 123869 171731 128968
rect 174966 123868 175310 128968
rect 176258 126840 176602 128968
rect 176258 126616 177386 126840
rect 178828 126774 179080 128968
rect 184037 126616 184289 128968
rect 176258 123868 176602 126616
rect 176985 125793 177364 125832
rect 176985 125646 177083 125793
rect 177255 125646 177364 125793
rect 176985 125608 177364 125646
rect 184119 125799 185113 125832
rect 184119 125652 184851 125799
rect 185023 125652 185113 125799
rect 184119 125608 185113 125652
rect 187622 123868 187966 128968
rect 188914 123868 189258 128968
rect 190371 123869 190715 128968
rect 193950 123868 194294 128968
rect 195242 123868 195586 128968
rect 196699 123869 197043 128968
rect 200278 123868 200622 128968
rect 201570 123868 201914 128968
rect 203027 128281 203371 128968
rect 204874 128545 205208 128968
rect 206612 128496 206946 128968
rect 208684 128468 209018 128968
rect 203027 128050 203102 128281
rect 203336 128050 203371 128281
rect 203027 126688 203371 128050
rect 215880 127533 217280 131263
rect 213318 127491 217289 127533
rect 213318 127238 213379 127491
rect 213645 127238 217289 127491
rect 213318 127198 217289 127238
rect 203027 126457 203089 126688
rect 203323 126457 203371 126688
rect 203027 125176 203371 126457
rect 215880 126044 217280 127198
rect 213309 125992 217280 126044
rect 213309 125739 213373 125992
rect 213639 125739 217280 125992
rect 213309 125709 217280 125739
rect 203027 124945 203067 125176
rect 203301 124945 203371 125176
rect 203027 123869 203371 124945
rect 215880 124267 217280 125709
rect 213302 124228 217280 124267
rect 213302 123975 213387 124228
rect 213653 123975 217280 124228
rect 213302 123932 217280 123975
rect 215880 121650 217280 123932
rect 152600 121557 162158 121650
rect 152600 121389 161759 121557
rect 161928 121389 162158 121557
rect 152600 121304 162158 121389
rect 206026 121304 217280 121650
rect 152600 120522 154000 121304
rect 206606 120960 206950 121062
rect 206606 120792 206696 120960
rect 206864 120792 206950 120960
rect 152600 120427 162158 120522
rect 152600 120259 161777 120427
rect 161946 120259 162158 120427
rect 206606 120284 206950 120792
rect 207255 120284 207599 121304
rect 207898 120960 208242 121062
rect 207898 120792 207984 120960
rect 208152 120792 208242 120960
rect 207898 120284 208242 120792
rect 208625 120277 208969 121304
rect 209355 120960 209699 121063
rect 209355 120792 209440 120960
rect 209608 120792 209699 120960
rect 209355 120285 209699 120792
rect 210080 120269 210424 121304
rect 152600 120176 162158 120259
rect 152600 118065 154000 120176
rect 215880 118066 217280 121304
rect 152600 117975 162158 118065
rect 152600 117807 161822 117975
rect 161991 117807 162158 117975
rect 152600 117719 162158 117807
rect 212240 117984 217280 118066
rect 212240 117816 212368 117984
rect 212537 117816 217280 117984
rect 212240 117720 217280 117816
rect 152600 116938 154000 117719
rect 215880 116938 217280 117720
rect 152600 116837 162158 116938
rect 152600 116669 161835 116837
rect 162004 116669 162158 116837
rect 152600 116592 162158 116669
rect 212240 116822 217280 116938
rect 212240 116654 212349 116822
rect 212518 116654 217280 116822
rect 212240 116592 217280 116654
rect 152600 114481 154000 116592
rect 215880 114482 217280 116592
rect 152600 114405 162158 114481
rect 152600 114237 161880 114405
rect 162049 114237 162158 114405
rect 152600 114135 162158 114237
rect 212240 114380 217280 114482
rect 212240 114212 212326 114380
rect 212495 114212 217280 114380
rect 212240 114136 217280 114212
rect 152600 113352 154000 114135
rect 215880 113354 217280 114136
rect 152600 113240 162158 113352
rect 152600 113072 161867 113240
rect 162036 113072 162158 113240
rect 152600 113006 162158 113072
rect 212240 113264 217280 113354
rect 212240 113096 212352 113264
rect 212521 113096 217280 113264
rect 212240 113008 217280 113096
rect 152600 105486 154000 113006
rect 158592 112504 158816 113006
rect 215880 110898 217280 113008
rect 212240 110802 217280 110898
rect 212240 110634 212326 110802
rect 212495 110634 217280 110802
rect 212240 110552 217280 110634
rect 215880 109770 217280 110552
rect 212240 109667 217280 109770
rect 212240 109499 212326 109667
rect 212495 109499 217280 109667
rect 212240 109424 217280 109499
rect 215880 107314 217280 109424
rect 212240 107183 217280 107314
rect 212240 107015 212355 107183
rect 212524 107015 217280 107183
rect 212240 106968 217280 107015
rect 215880 106186 217280 106968
rect 212240 106066 217280 106186
rect 212240 105898 212323 106066
rect 212492 105898 217280 106066
rect 212240 105840 217280 105898
rect 158592 105486 158816 105735
rect 152600 105140 158816 105486
rect 152600 103727 154000 105140
rect 215880 103730 217280 105840
rect 152600 103647 162158 103727
rect 152600 103479 161804 103647
rect 161973 103479 162158 103647
rect 152600 103381 162158 103479
rect 212240 103611 217280 103730
rect 212240 103443 212346 103611
rect 212515 103443 217280 103611
rect 212240 103384 217280 103443
rect 152600 102602 154000 103381
rect 215880 102602 217280 103384
rect 152600 102488 162158 102602
rect 152600 102320 161837 102488
rect 162006 102320 162158 102488
rect 152600 102256 162158 102320
rect 212240 102498 217280 102602
rect 212240 102330 212336 102498
rect 212505 102330 217280 102498
rect 212240 102256 217280 102330
rect 152600 100145 154000 102256
rect 215880 100146 217280 102256
rect 152600 100056 162158 100145
rect 152600 99888 161822 100056
rect 161991 99888 162158 100056
rect 152600 99799 162158 99888
rect 212240 100040 217280 100146
rect 212240 99872 212342 100040
rect 212511 99872 217280 100040
rect 212240 99800 217280 99872
rect 152600 99025 154000 99799
rect 152600 98912 162158 99025
rect 215880 99018 217280 99800
rect 152600 98744 161870 98912
rect 162039 98744 162158 98912
rect 152600 98679 162158 98744
rect 212240 98911 217280 99018
rect 212240 98743 212342 98911
rect 212511 98743 217280 98911
rect 152600 96561 154000 98679
rect 212240 98672 217280 98743
rect 215880 96562 217280 98672
rect 152600 96477 162158 96561
rect 152600 96309 161808 96477
rect 161977 96309 162158 96477
rect 152600 96215 162158 96309
rect 212240 96475 217280 96562
rect 212240 96307 212349 96475
rect 212518 96307 217280 96475
rect 212240 96216 217280 96307
rect 152600 95434 154000 96215
rect 215880 95434 217280 96216
rect 152600 95306 162158 95434
rect 152600 95138 161780 95306
rect 161949 95138 162158 95306
rect 152600 95088 162158 95138
rect 212240 95365 217280 95434
rect 212240 95197 212363 95365
rect 212532 95197 217280 95365
rect 212240 95088 217280 95197
rect 152600 91557 154000 95088
rect 162310 94248 162654 94595
rect 163602 94248 163946 94590
rect 165059 94248 165404 94626
rect 168639 94248 168984 94612
rect 169929 94248 170274 94620
rect 171387 94248 171732 94626
rect 174966 94248 175311 94605
rect 176258 94248 176603 94603
rect 177715 94248 178060 94605
rect 181294 94248 181639 94611
rect 182586 94248 182931 94617
rect 184043 94248 184388 94589
rect 187622 94248 187967 94624
rect 188914 94248 189259 94600
rect 190371 94248 190716 94609
rect 193949 94248 194294 94618
rect 195242 94248 195587 94612
rect 196698 94248 197043 94619
rect 200277 94248 200622 94608
rect 201570 94248 201915 94608
rect 203026 94248 203371 94615
rect 206605 94248 206950 94613
rect 207897 94248 208242 94616
rect 209355 94248 209700 94611
rect 154952 93960 215320 94248
rect 154952 93851 214245 93960
rect 154952 93096 155263 93851
rect 156044 93205 214245 93851
rect 215026 93205 215320 93960
rect 156044 93096 215320 93205
rect 154952 92848 215320 93096
rect 152600 90802 152887 91557
rect 153668 90802 154000 91557
rect 152600 90552 154000 90802
rect 215880 91557 217280 95088
rect 215880 90802 216239 91557
rect 217020 90802 217280 91557
rect 215880 90552 217280 90802
<< via3 >>
rect 152901 131298 153682 132053
rect 216237 131263 217018 132018
rect 155290 129236 156071 129991
rect 214286 129264 215067 130019
rect 177083 125646 177255 125793
rect 184851 125652 185023 125799
rect 203102 128050 203336 128281
rect 213379 127238 213645 127491
rect 203089 126457 203323 126688
rect 213373 125739 213639 125992
rect 203067 124945 203301 125176
rect 213387 123975 213653 124228
rect 163072 123312 163184 123424
rect 164436 123312 164548 123424
rect 165892 123312 166004 123424
rect 169400 123312 169512 123424
rect 170768 123312 170880 123424
rect 172230 123312 172342 123424
rect 175728 123312 175840 123424
rect 177096 123312 177208 123424
rect 178553 123312 178665 123424
rect 182056 123312 182168 123424
rect 183426 123312 183538 123424
rect 184884 123312 184996 123424
rect 188384 123312 188496 123424
rect 189757 123312 189869 123424
rect 191208 123312 191320 123424
rect 194712 123312 194824 123424
rect 196083 123312 196195 123424
rect 197540 123312 197652 123424
rect 201040 123312 201152 123424
rect 202414 123312 202526 123424
rect 161759 121389 161928 121557
rect 206696 120792 206864 120960
rect 161777 120259 161946 120427
rect 207984 120792 208152 120960
rect 209440 120792 209608 120960
rect 161822 117807 161991 117975
rect 212368 117816 212537 117984
rect 161835 116669 162004 116837
rect 212349 116654 212518 116822
rect 161880 114237 162049 114405
rect 212326 114212 212495 114380
rect 161867 113072 162036 113240
rect 212352 113096 212521 113264
rect 157648 112343 157753 112447
rect 157640 112001 157752 112057
rect 212326 110634 212495 110802
rect 212326 109499 212495 109667
rect 157640 108473 157752 108529
rect 212355 107015 212524 107183
rect 157640 106625 157752 106681
rect 212323 105898 212492 106066
rect 161804 103479 161973 103647
rect 212346 103443 212515 103611
rect 161837 102320 162006 102488
rect 212336 102330 212505 102498
rect 161822 99888 161991 100056
rect 212342 99872 212511 100040
rect 161870 98744 162039 98912
rect 212342 98743 212511 98911
rect 161808 96309 161977 96477
rect 212349 96307 212518 96475
rect 161780 95138 161949 95306
rect 212363 95197 212532 95365
rect 155263 93096 156044 93851
rect 214245 93205 215026 93960
rect 152887 90802 153668 91557
rect 216239 90802 217020 91557
<< metal4 >>
rect 152600 132053 217282 132384
rect 152600 131298 152901 132053
rect 153682 132018 217282 132053
rect 153682 131298 216237 132018
rect 152600 131263 216237 131298
rect 217018 131263 217282 132018
rect 152600 130984 217282 131263
rect 154952 129991 156352 130368
rect 154952 129236 155290 129991
rect 156071 129236 156352 129991
rect 154952 122290 156352 129236
rect 162959 123424 163304 130984
rect 162959 123312 163072 123424
rect 163184 123312 163304 123424
rect 162959 123256 163304 123312
rect 164329 123424 164674 130984
rect 164329 123312 164436 123424
rect 164548 123312 164674 123424
rect 164329 123256 164674 123312
rect 165784 123424 166129 130984
rect 165784 123312 165892 123424
rect 166004 123312 166129 123424
rect 165784 123256 166129 123312
rect 169287 123424 169632 130984
rect 169287 123312 169400 123424
rect 169512 123312 169632 123424
rect 169287 123256 169632 123312
rect 170657 123424 171002 130984
rect 170657 123312 170768 123424
rect 170880 123312 171002 123424
rect 170657 123256 171002 123312
rect 172112 123424 172457 130984
rect 172112 123312 172230 123424
rect 172342 123312 172457 123424
rect 172112 123256 172457 123312
rect 175616 123424 175961 130984
rect 175616 123312 175728 123424
rect 175840 123312 175961 123424
rect 175616 123256 175961 123312
rect 176985 125793 177330 130984
rect 176985 125646 177083 125793
rect 177255 125646 177330 125793
rect 176985 123424 177330 125646
rect 176985 123312 177096 123424
rect 177208 123312 177330 123424
rect 176985 123256 177330 123312
rect 178440 123424 178785 130984
rect 178440 123312 178553 123424
rect 178665 123312 178785 123424
rect 178440 123256 178785 123312
rect 181943 123424 182288 130984
rect 181943 123312 182056 123424
rect 182168 123312 182288 123424
rect 181943 123256 182288 123312
rect 183313 123424 183658 130984
rect 183313 123312 183426 123424
rect 183538 123312 183658 123424
rect 183313 123255 183658 123312
rect 184767 125799 185112 130984
rect 184767 125652 184851 125799
rect 185023 125652 185112 125799
rect 184767 123424 185112 125652
rect 184767 123312 184884 123424
rect 184996 123312 185112 123424
rect 184767 123255 185112 123312
rect 188271 123424 188616 130984
rect 188271 123312 188384 123424
rect 188496 123312 188616 123424
rect 188271 123256 188616 123312
rect 189641 123424 189986 130984
rect 189641 123312 189757 123424
rect 189869 123312 189986 123424
rect 189641 123256 189986 123312
rect 191096 123424 191441 130984
rect 191096 123312 191208 123424
rect 191320 123312 191441 123424
rect 191096 123256 191441 123312
rect 194599 123424 194944 130984
rect 194599 123312 194712 123424
rect 194824 123312 194944 123424
rect 194599 123256 194944 123312
rect 195969 123424 196314 130984
rect 195969 123312 196083 123424
rect 196195 123312 196314 123424
rect 195969 123256 196314 123312
rect 197424 123424 197769 130984
rect 197424 123312 197540 123424
rect 197652 123312 197769 123424
rect 197424 123256 197769 123312
rect 200927 123424 201272 130984
rect 200927 123312 201040 123424
rect 201152 123312 201272 123424
rect 200927 123256 201272 123312
rect 202297 127536 202642 130984
rect 213920 130019 215320 130368
rect 213920 129264 214286 130019
rect 215067 129264 215320 130019
rect 213920 128329 215320 129264
rect 203024 128281 204471 128328
rect 203024 128050 203102 128281
rect 203336 128050 204471 128281
rect 203024 127995 204471 128050
rect 213750 127994 215320 128329
rect 202297 127203 204080 127536
rect 202297 126042 202642 127203
rect 213920 126744 215320 127994
rect 203028 126688 204475 126741
rect 203028 126457 203089 126688
rect 203323 126457 204475 126688
rect 203028 126408 204475 126457
rect 213769 126409 215320 126744
rect 202297 125709 204059 126042
rect 202297 124268 202642 125709
rect 213920 125248 215320 126409
rect 203025 125176 204472 125247
rect 203025 124945 203067 125176
rect 203301 124945 204472 125176
rect 203025 124914 204472 124945
rect 213810 124913 215320 125248
rect 202297 123935 204074 124268
rect 202297 123424 202642 123935
rect 202297 123312 202414 123424
rect 202526 123312 202642 123424
rect 202297 123256 202642 123312
rect 154952 121943 161075 122290
rect 213920 122289 215320 124913
rect 206451 121944 215320 122289
rect 154952 121063 156352 121943
rect 154952 120716 161067 121063
rect 213920 121062 215320 121944
rect 206470 120960 215320 121062
rect 206470 120792 206696 120960
rect 206864 120792 207984 120960
rect 208152 120792 209440 120960
rect 209608 120792 215320 120960
rect 206470 120717 215320 120792
rect 154952 118706 156352 120716
rect 154952 118359 161075 118706
rect 213920 118705 215320 120717
rect 212778 118360 215320 118705
rect 154952 117479 156352 118359
rect 154952 117132 161067 117479
rect 213920 117478 215320 118360
rect 212798 117133 215320 117478
rect 154952 115122 156352 117132
rect 154952 114775 161075 115122
rect 213920 115121 215320 117133
rect 212779 114776 215320 115121
rect 154952 113895 156352 114775
rect 154952 113548 161067 113895
rect 213920 113894 215320 114776
rect 212798 113549 215320 113894
rect 154952 112128 156352 113548
rect 157584 112447 157808 113548
rect 157584 112343 157648 112447
rect 157753 112343 157808 112447
rect 157584 112294 157808 112343
rect 154952 112057 157835 112128
rect 154952 112001 157640 112057
rect 157752 112001 157835 112057
rect 154952 111948 157835 112001
rect 154952 111538 156352 111948
rect 154952 111191 161075 111538
rect 213920 111537 215320 113549
rect 212779 111192 215320 111537
rect 154952 110311 156352 111191
rect 213920 110311 215320 111192
rect 154952 109964 161067 110311
rect 213684 110310 215320 110311
rect 212798 109966 215320 110310
rect 212798 109965 213696 109966
rect 154952 108618 156352 109964
rect 154952 108529 158003 108618
rect 154952 108473 157640 108529
rect 157752 108473 158003 108529
rect 154952 108385 158003 108473
rect 154952 107953 156352 108385
rect 213920 107953 215320 109966
rect 154952 107606 161075 107953
rect 212779 107608 215320 107953
rect 154952 106727 156352 107606
rect 154952 106681 161067 106727
rect 213920 106726 215320 107608
rect 154952 106625 157640 106681
rect 157752 106625 161067 106681
rect 154952 106380 161067 106625
rect 212798 106381 215320 106726
rect 154952 104370 156352 106380
rect 154952 104023 161075 104370
rect 213920 104369 215320 106381
rect 212779 104024 215320 104369
rect 154952 103143 156352 104023
rect 154952 102796 161067 103143
rect 213920 103142 215320 104024
rect 212798 102797 215320 103142
rect 154952 100786 156352 102796
rect 154952 100439 161075 100786
rect 213920 100785 215320 102797
rect 212779 100440 215320 100785
rect 154952 99559 156352 100439
rect 154952 99212 161067 99559
rect 213920 99558 215320 100440
rect 212798 99213 215320 99558
rect 154952 97202 156352 99212
rect 154952 96855 161075 97202
rect 213920 97201 215320 99213
rect 212779 96856 215320 97201
rect 154952 95975 156352 96855
rect 154952 95628 161067 95975
rect 213920 95974 215320 96856
rect 212798 95629 215320 95974
rect 154952 93851 156352 95628
rect 154952 93096 155263 93851
rect 156044 93096 156352 93851
rect 154952 92848 156352 93096
rect 162959 91952 163303 95088
rect 164329 91952 164673 95088
rect 165784 91952 166128 95088
rect 169287 91952 169631 95088
rect 170657 91952 171001 95088
rect 172112 91952 172456 95088
rect 175615 91952 175959 95088
rect 176985 91952 177329 95088
rect 178440 91952 178784 95088
rect 181943 91952 182287 95088
rect 183313 91952 183657 95088
rect 184768 91952 185112 95088
rect 188271 91952 188615 95088
rect 189641 91952 189985 95089
rect 191096 91952 191440 95088
rect 194599 91952 194943 95088
rect 195969 91952 196313 95088
rect 197424 91952 197768 95088
rect 200927 91952 201271 95088
rect 202297 91952 202641 95088
rect 203752 91952 204096 95088
rect 207255 91952 207599 95088
rect 208625 91952 208969 95088
rect 210080 91952 210424 95088
rect 213920 93960 215320 95629
rect 213920 93205 214245 93960
rect 215026 93205 215320 93960
rect 213920 92848 215320 93205
rect 152600 91557 217280 91952
rect 152600 90802 152887 91557
rect 153668 90802 216239 91557
rect 217020 90802 217280 91557
rect 152600 90552 217280 90802
use 4MSB_weighted_binary  4MSB_weighted_binary_0
timestamp 1758278152
transform 1 0 202104 0 1 126824
box 1838 -3064 11724 1721
use 6MSB_MATRIX  6MSB_MATRIX_0
timestamp 1758622385
transform 1 0 120680 0 1 81760
box 40152 12656 92904 42109
use thermo_decoder  thermo_decoder_0
timestamp 1757908133
transform 1 0 156128 0 1 106065
box 336 -337 3920 6440
use thermo_decoder  thermo_decoder_1
timestamp 1757908133
transform 0 1 177689 -1 0 128296
box 336 -337 3920 6440
<< labels >>
flabel metal2 205637 132386 205790 132532 1 FreeSans 4800 0 0 0 X1
port 1 n
flabel metal2 203738 132396 203891 132542 1 FreeSans 4800 0 0 0 X2
port 2 n
flabel metal2 202337 132396 202490 132542 1 FreeSans 4800 0 0 0 X3
port 3 n
flabel metal2 200544 132390 200697 132536 1 FreeSans 4800 0 0 0 X4
port 4 n
flabel metal2 184808 132398 184961 132544 1 FreeSans 4800 0 0 0 X5
port 5 n
flabel metal1 180609 132391 180762 132537 1 FreeSans 4800 0 0 0 X6
port 6 n
flabel metal1 176912 132394 177065 132540 1 FreeSans 4800 0 0 0 X7
port 7 n
flabel metal1 159664 132397 159817 132543 1 FreeSans 4800 0 0 0 X10
port 10 n
flabel metal2 156805 132395 156958 132541 1 FreeSans 4800 0 0 0 X8
port 8 n
flabel metal1 156473 131546 156626 131692 1 FreeSans 4800 0 0 0 X9
port 9 n
flabel metal1 188670 132404 188821 132541 1 FreeSans 4800 0 0 0 CLK
port 11 n
flabel metal1 212381 132390 212666 132522 1 FreeSans 4800 0 0 0 OUTP
port 12 n
flabel metal1 212833 131508 213118 131640 1 FreeSans 4800 0 0 0 OUTN
port 13 n
flabel metal1 213276 130712 213561 130844 1 FreeSans 4800 0 0 0 VBIAS
port 14 n
flabel metal3 154952 128968 215320 130368 1 FreeSans 8000 0 0 0 VDD
port 15 n
flabel metal4 213920 92848 215320 130368 1 FreeSans 8000 0 0 0 VDD
port 15 n
flabel metal3 154952 92848 215320 94248 1 FreeSans 8000 0 0 0 VDD
port 15 n
flabel metal4 154952 92848 156352 130368 1 FreeSans 8000 0 0 0 VDD
port 15 n
flabel metal3 215880 90552 217280 132384 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel metal4 152600 90552 217280 91952 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel metal3 152600 90552 154000 132384 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel metal4 152600 130984 217282 132384 1 FreeSans 8000 0 0 0 VSS
port 16 n
<< end >>
