* SPICE3 file created from CS_Switch_16x.ext - technology: gf180mcuD

.subckt CS_Switch_16x INP INN OUTP OUTN VBIAS VSS VPW
X0 a_1640_n12# VBIAS a_1304_n132# VPW nfet_03v3 ad=0.1357p pd=1.08u as=0.2264p ps=2.1u w=0.56u l=0.28u
X1 VSS VBIAS a_1640_n12# VPW nfet_03v3 ad=0.2358p pd=2.18u as=0.1357p ps=1.08u w=0.62u l=0.3u
X2 VSS VBIAS a_1640_n192# VPW nfet_03v3 ad=0.2358p pd=2.18u as=0.1357p ps=1.08u w=0.62u l=0.3u
X3 OUTN INN a_1304_n132# VPW nfet_03v3 ad=0.234p pd=2.14u as=0.218p ps=1.66u w=0.6u l=0.3u
X4 a_1304_n132# INP OUTP VPW nfet_03v3 ad=0.218p pd=1.66u as=0.234p ps=2.14u w=0.6u l=0.3u
X5 a_1640_n192# VBIAS a_1304_n132# VPW nfet_03v3 ad=0.1357p pd=1.08u as=0.2264p ps=2.1u w=0.56u l=0.28u
C0 INP INN 0.058006f
C1 INP VBIAS 0.001437f
C2 INN VBIAS 0.001551f
C3 VSS a_1640_n192# 0.007182f
C4 INN a_1640_n12# 0.001013f
C5 OUTN INP 3.49e-19
C6 OUTP INP 0.007401f
C7 OUTN INN 0.007874f
C8 OUTP INN 3.2e-19
C9 VBIAS a_1640_n12# 0.00422f
C10 OUTN VBIAS 0.019262f
C11 INP a_1304_n132# 0.00715f
C12 OUTP VBIAS 0.00181f
C13 INN a_1304_n132# 0.00715f
C14 OUTN OUTP 0.002923f
C15 a_1304_n132# VBIAS 0.007442f
C16 INP VSS 0.038477f
C17 VSS INN 7.92e-19
C18 a_1304_n132# a_1640_n12# 2.3e-19
C19 OUTN a_1304_n132# 0.04805f
C20 OUTP a_1304_n132# 0.046263f
C21 VSS VBIAS 0.045797f
C22 INP a_1640_n192# 0.001013f
C23 VSS a_1640_n12# 0.002225f
C24 OUTN VSS 1.82e-19
C25 OUTP VSS 0.159563f
C26 VBIAS a_1640_n192# 0.002733f
C27 VSS a_1304_n132# 0.034263f
C28 a_1304_n132# a_1640_n192# 2.3e-19
C29 OUTP VPW 0.028916f
C30 INP VPW 0.229072f
C31 VSS VPW 0.428197f
C32 INN VPW 0.246194f
C33 OUTN VPW 0.056853f
C34 VBIAS VPW 0.504283f
C35 a_1304_n132# VPW 0.04863f
.ends

