magic
tech gf180mcuD
magscale 1 10
timestamp 1754627642
<< isosubstrate >>
rect 518 1526 1757 2149
<< pwell >>
rect 518 1526 1757 2149
<< nmos >>
rect 644 1918 700 1962
rect 1040 1918 1096 1962
rect 1180 1918 1236 1962
rect 644 1708 700 1770
rect 894 1708 954 1770
rect 1576 1918 1632 1962
rect 1040 1710 1096 1766
rect 1180 1710 1236 1766
rect 1320 1708 1380 1770
rect 1576 1708 1632 1770
<< ndiff >>
rect 940 1963 1020 1980
rect 560 1918 644 1962
rect 700 1918 746 1962
rect 940 1917 957 1963
rect 1003 1962 1020 1963
rect 1256 1963 1336 1980
rect 1256 1962 1273 1963
rect 1003 1918 1040 1962
rect 1096 1918 1180 1962
rect 1236 1918 1273 1962
rect 1003 1917 1020 1918
rect 940 1900 1020 1917
rect 802 1770 874 1780
rect 598 1708 644 1770
rect 700 1708 746 1770
rect 802 1767 894 1770
rect 802 1721 815 1767
rect 861 1721 894 1767
rect 802 1708 894 1721
rect 954 1766 1004 1770
rect 1116 1766 1160 1918
rect 1256 1917 1273 1918
rect 1319 1917 1336 1963
rect 1530 1918 1576 1962
rect 1632 1918 1716 1962
rect 1256 1900 1336 1917
rect 1402 1770 1474 1780
rect 1272 1766 1320 1770
rect 954 1710 1040 1766
rect 1096 1710 1180 1766
rect 1236 1710 1320 1766
rect 954 1708 1020 1710
rect 976 1634 1020 1708
rect 1256 1708 1320 1710
rect 1380 1767 1474 1770
rect 1380 1721 1415 1767
rect 1461 1721 1474 1767
rect 1380 1708 1474 1721
rect 1530 1708 1576 1770
rect 1632 1708 1678 1770
rect 1256 1634 1300 1708
rect 976 1590 1300 1634
<< ndiffc >>
rect 957 1917 1003 1963
rect 815 1721 861 1767
rect 1273 1917 1319 1963
rect 1415 1721 1461 1767
<< polysilicon >>
rect 1028 2087 1108 2104
rect 1028 2041 1045 2087
rect 1091 2041 1108 2087
rect 1028 2024 1108 2041
rect 1168 2087 1248 2104
rect 1168 2041 1185 2087
rect 1231 2041 1248 2087
rect 1168 2024 1248 2041
rect 644 1962 700 2008
rect 644 1770 700 1918
rect 1040 1962 1096 2024
rect 1180 1962 1236 2024
rect 816 1885 896 1902
rect 816 1839 833 1885
rect 879 1858 896 1885
rect 1040 1874 1096 1918
rect 879 1839 930 1858
rect 816 1826 930 1839
rect 816 1822 1096 1826
rect 894 1790 1096 1822
rect 894 1770 954 1790
rect 1040 1766 1096 1790
rect 1180 1874 1236 1918
rect 1576 1962 1632 2008
rect 1380 1885 1460 1902
rect 1380 1858 1397 1885
rect 1344 1839 1397 1858
rect 1443 1839 1460 1885
rect 1344 1826 1460 1839
rect 1180 1822 1460 1826
rect 1180 1790 1380 1822
rect 1180 1766 1236 1790
rect 1320 1770 1380 1790
rect 1576 1770 1632 1918
rect 644 1664 700 1708
rect 636 1651 708 1664
rect 894 1662 954 1708
rect 636 1605 649 1651
rect 695 1605 708 1651
rect 636 1592 708 1605
rect 1040 1690 1096 1710
rect 1180 1690 1236 1710
rect 1040 1654 1236 1690
rect 1320 1662 1380 1708
rect 1576 1662 1632 1708
rect 1568 1649 1640 1662
rect 1568 1603 1581 1649
rect 1627 1603 1640 1649
rect 1568 1590 1640 1603
<< polycontact >>
rect 1045 2041 1091 2087
rect 1185 2041 1231 2087
rect 833 1839 879 1885
rect 1397 1839 1443 1885
rect 649 1605 695 1651
rect 1581 1603 1627 1649
<< metal1 >>
rect 1030 2087 1106 2102
rect 1030 2041 1045 2087
rect 1091 2041 1106 2087
rect 1030 2026 1106 2041
rect 1170 2087 1246 2102
rect 1170 2041 1185 2087
rect 1231 2041 1246 2087
rect 1170 2026 1246 2041
rect 942 1963 1018 1978
rect 942 1917 957 1963
rect 1003 1917 1018 1963
rect 942 1902 1018 1917
rect 1258 1963 1334 1978
rect 1258 1917 1273 1963
rect 1319 1917 1334 1963
rect 1258 1902 1334 1917
rect 818 1885 894 1900
rect 818 1839 833 1885
rect 879 1839 894 1885
rect 818 1824 894 1839
rect 1382 1885 1458 1900
rect 1382 1839 1397 1885
rect 1443 1839 1458 1885
rect 1382 1824 1458 1839
rect 815 1767 861 1778
rect 815 1686 861 1721
rect 1415 1767 1461 1778
rect 1415 1686 1461 1721
rect 596 1651 1690 1686
rect 596 1605 649 1651
rect 695 1649 1690 1651
rect 695 1605 1581 1649
rect 596 1603 1581 1605
rect 1627 1603 1690 1649
rect 596 1566 1690 1603
<< labels >>
flabel metal1 1030 2026 1106 2102 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 1170 2026 1246 2102 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 942 1902 1018 1978 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 1258 1902 1334 1978 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 818 1824 894 1900 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 1382 1824 1458 1900 1 FreeSans 400 0 0 0 VBIAS
port 6 nsew power bidirectional
flabel metal1 788 1566 1481 1686 1 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional
flabel pwell 1436 1550 1515 1696 1 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
<< end >>
