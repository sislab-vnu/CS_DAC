magic
tech gf180mcuD
magscale 1 10
timestamp 1755843645
<< nwell >>
rect 1227 249 1452 253
rect 1228 167 1444 249
rect 1227 -230 1452 167
rect 2512 -261 2830 253
<< pwell >>
rect 1279 253 1497 691
rect 2586 253 2881 691
<< psubdiff >>
rect 1253 636 1421 660
rect 1253 577 1294 636
rect 1382 577 1421 636
rect 1253 552 1421 577
rect 2615 627 2767 651
rect 2615 566 2643 627
rect 2738 566 2767 627
rect 2615 550 2767 566
rect 77 -1056 190 -1029
rect 77 -1123 98 -1056
rect 167 -1123 190 -1056
rect 77 -1138 190 -1123
<< nsubdiff >>
rect 87 -226 212 -195
rect 87 -293 109 -226
rect 189 -293 212 -226
rect 87 -320 212 -293
rect 3418 -212 3534 -192
rect 3418 -279 3435 -212
rect 3515 -279 3534 -212
rect 3418 -303 3534 -279
<< psubdiffcont >>
rect 1294 577 1382 636
rect 2643 566 2738 627
rect 98 -1123 167 -1056
<< nsubdiffcont >>
rect 109 -293 189 -226
rect 3435 -279 3515 -212
<< metal1 >>
rect 1193 636 1516 665
rect 1193 577 1294 636
rect 1382 577 1516 636
rect 1193 545 1516 577
rect 2519 627 3164 665
rect 2519 566 2643 627
rect 2738 566 3164 627
rect 2519 545 3164 566
rect 3410 69 4364 133
rect 1192 -240 1544 -119
rect 2508 -239 2882 -119
rect 2508 -240 2860 -239
rect 3661 -554 4190 -493
rect 4300 -495 4364 69
rect 3661 -617 3722 -554
rect 3356 -678 3722 -617
rect 3539 -1143 3797 -1023
<< via1 >>
rect 3043 198 3287 252
rect 1766 -61 1820 97
rect 1004 -809 1056 -576
rect 3176 -590 3324 -526
<< metal2 >>
rect 3000 252 3304 264
rect 3000 198 3043 252
rect 3287 198 3304 252
rect 3000 181 3304 198
rect 1758 97 1830 133
rect 1758 -38 1766 97
rect 988 -61 1766 -38
rect 1820 -61 1830 97
rect 988 -119 1830 -61
rect 988 -576 1069 -119
rect 988 -809 1004 -576
rect 1056 -809 1069 -576
rect 3140 -488 3219 181
rect 3140 -526 3356 -488
rect 3140 -590 3176 -526
rect 3324 -590 3356 -526
rect 3140 -617 3356 -590
rect 988 -841 1069 -809
use CS_Switch_16x2  CS_Switch_16x2_0
timestamp 1755760707
transform 1 0 4009 0 1 -1833
box -377 631 825 1384
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 74 0 1 -1083
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2874 0 -1 605
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  gf180mcu_fd_sc_mcu7t5v0__nand2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 1514 0 -1 605
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 74 0 -1 605
box -86 -86 1206 870
<< end >>
