* NGSPICE file created from CS_Switch_2x2.ext - technology: gf180mcuD

.subckt CS_Switch_2x2 INP INN OUTP OUTN VBIAS VSS
X0 a_336_n248# VBIAS a_32_n20# VSS nfet_03v3 ad=0.2728p pd=1.905u as=0.1516p ps=1.64u w=0.22u l=0.28u
X1 OUTN INN a_32_n20# VSS nfet_03v3 ad=0.182p pd=1.8u as=0.102p ps=1u w=0.22u l=0.28u
X2 a_32_n20# INP OUTP VSS nfet_03v3 ad=0.102p pd=1u as=0.102p ps=1u w=0.22u l=0.28u
X3 OUTP VSS a_n246_n20# VSS nfet_03v3 ad=0.102p pd=1u as=50.6f ps=0.9u w=0.22u l=0.28u
X4 a_336_n248# VBIAS VSS VSS nfet_03v3 ad=0.2728p pd=1.905u as=0.132p ps=1.04u w=0.44u l=1.8u
X5 a_652_n20# VSS a_336_n248# VSS nfet_03v3 ad=50.6f pd=0.9u as=0.2728p ps=1.905u w=0.22u l=0.28u
X6 a_652_n248# VSS a_336_n248# VSS nfet_03v3 ad=0.1012p pd=1.34u as=0.2728p ps=1.905u w=0.44u l=0.28u
X7 VSS VSS a_n246_n248# VSS nfet_03v3 ad=0.132p pd=1.04u as=0.1012p ps=1.34u w=0.44u l=0.28u
C0 INN OUTP 7.31e-20
C1 OUTN VBIAS 0.001721f
C2 a_n246_n20# OUTP 7.78e-19
C3 a_336_n248# VBIAS 0.001759f
C4 OUTN a_32_n20# 0.163167f
C5 INP OUTN 7.31e-20
C6 a_32_n20# a_336_n248# 0.004758f
C7 a_32_n20# VBIAS 0.049088f
C8 INP VBIAS 0.019794f
C9 INP a_32_n20# 0.003036f
C10 OUTN OUTP 6.13e-19
C11 INN OUTN 0.003859f
C12 a_32_n20# OUTP 0.028781f
C13 INP OUTP 0.003859f
C14 INN VBIAS 0.041085f
C15 INN a_32_n20# 0.029571f
C16 INN INP 0.055413f
C17 OUTN VSS 0.018799f
C18 OUTP VSS 0.059535f
C19 VBIAS VSS 0.903508f
C20 INN VSS 0.178433f
C21 INP VSS 0.211357f
C22 a_652_n248# VSS 0.001884f
C23 a_n246_n248# VSS 0.00298f
C24 a_652_n20# VSS 4.96e-19
C25 a_336_n248# VSS 0.014638f
C26 a_n246_n20# VSS 4.96e-19
C27 a_32_n20# VSS 0.217029f
.ends

