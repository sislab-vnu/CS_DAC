magic
tech gf180mcuD
magscale 1 10
timestamp 1754365189
<< pwell >>
rect -376 -1440 992 -520
<< nmos >>
rect -169 -827 -113 -783
rect 59 -827 115 -783
rect 448 -849 808 -759
rect -170 -1050 -114 -1006
rect 58 -1050 114 -1006
rect 448 -1073 808 -983
<< ndiff >>
rect -295 -783 -215 -765
rect -67 -783 13 -765
rect 402 -765 448 -759
rect 161 -780 241 -765
rect 161 -783 179 -780
rect -295 -784 -169 -783
rect -295 -830 -279 -784
rect -233 -827 -169 -784
rect -113 -827 -50 -783
rect -233 -830 -215 -827
rect -295 -845 -215 -830
rect -67 -829 -50 -827
rect -4 -827 59 -783
rect 115 -826 179 -783
rect 225 -826 241 -780
rect 115 -827 241 -826
rect -4 -829 13 -827
rect -67 -845 13 -829
rect 161 -845 241 -827
rect 322 -780 448 -765
rect 322 -826 340 -780
rect 386 -826 448 -780
rect 322 -845 448 -826
rect 402 -849 448 -845
rect 808 -763 854 -759
rect 808 -778 934 -763
rect 808 -824 872 -778
rect 918 -824 934 -778
rect 808 -843 934 -824
rect 808 -849 854 -843
rect -296 -1006 -216 -988
rect -68 -1004 12 -988
rect -68 -1006 -51 -1004
rect -296 -1007 -170 -1006
rect -296 -1053 -280 -1007
rect -234 -1050 -170 -1007
rect -114 -1050 -51 -1006
rect -5 -1006 12 -1004
rect 160 -1003 240 -988
rect 402 -989 448 -983
rect 160 -1006 178 -1003
rect -5 -1050 58 -1006
rect 114 -1049 178 -1006
rect 224 -1049 240 -1003
rect 114 -1050 240 -1049
rect -234 -1053 -216 -1050
rect -296 -1068 -216 -1053
rect -68 -1068 12 -1050
rect 160 -1068 240 -1050
rect 322 -1004 448 -989
rect 322 -1050 340 -1004
rect 386 -1050 448 -1004
rect 322 -1069 448 -1050
rect 402 -1073 448 -1069
rect 808 -988 854 -983
rect 808 -1003 934 -988
rect 808 -1049 872 -1003
rect 918 -1049 934 -1003
rect 808 -1068 934 -1049
rect 808 -1073 854 -1068
<< ndiffc >>
rect -279 -830 -233 -784
rect -50 -829 -4 -783
rect 179 -826 225 -780
rect 340 -826 386 -780
rect 872 -824 918 -778
rect -280 -1053 -234 -1007
rect -51 -1050 -5 -1004
rect 178 -1049 224 -1003
rect 340 -1050 386 -1004
rect 872 -1049 918 -1003
<< polysilicon >>
rect -180 -675 -100 -657
rect -180 -721 -163 -675
rect -117 -721 -100 -675
rect -180 -737 -100 -721
rect 48 -675 128 -657
rect 48 -721 65 -675
rect 111 -721 128 -675
rect 48 -737 128 -721
rect -169 -783 -113 -737
rect 59 -783 115 -737
rect 448 -759 808 -713
rect -169 -873 -113 -827
rect 59 -873 115 -827
rect 448 -896 808 -849
rect 448 -942 573 -896
rect 693 -942 808 -896
rect -170 -1006 -114 -960
rect 58 -1006 114 -960
rect 448 -983 808 -942
rect -170 -1098 -114 -1050
rect 58 -1098 114 -1050
rect 448 -1098 808 -1073
rect -170 -1134 808 -1098
rect 488 -1135 808 -1134
<< polycontact >>
rect -163 -721 -117 -675
rect 65 -721 111 -675
rect 573 -942 693 -896
<< metal1 >>
rect -284 -767 -228 -615
rect -169 -675 -110 -616
rect -169 -721 -163 -675
rect -117 -721 -110 -675
rect -169 -732 -110 -721
rect 55 -675 114 -616
rect 55 -721 65 -675
rect 111 -721 114 -675
rect 55 -732 114 -721
rect 174 -767 230 -612
rect -294 -784 -218 -767
rect -294 -830 -279 -784
rect -233 -830 -218 -784
rect -294 -843 -218 -830
rect -65 -783 11 -767
rect -65 -829 -50 -783
rect -4 -829 11 -783
rect -65 -843 11 -829
rect 164 -780 240 -767
rect 164 -826 179 -780
rect 225 -826 240 -780
rect 164 -843 240 -826
rect 325 -780 401 -767
rect 325 -826 340 -780
rect 386 -826 401 -780
rect 325 -843 401 -826
rect 857 -778 933 -765
rect 857 -824 872 -778
rect 918 -824 933 -778
rect 857 -841 933 -824
rect -51 -990 -4 -843
rect 340 -895 386 -843
rect 178 -941 386 -895
rect 505 -896 777 -884
rect 178 -990 224 -941
rect 505 -942 573 -896
rect 693 -942 777 -896
rect 505 -953 777 -942
rect 872 -990 918 -841
rect -295 -1007 -219 -990
rect -295 -1053 -280 -1007
rect -234 -1053 -219 -1007
rect -295 -1066 -219 -1053
rect -66 -1004 10 -990
rect -66 -1050 -51 -1004
rect -5 -1050 10 -1004
rect -66 -1066 10 -1050
rect 163 -1003 239 -990
rect 163 -1049 178 -1003
rect 224 -1049 239 -1003
rect 163 -1066 239 -1049
rect 325 -1004 401 -991
rect 325 -1050 340 -1004
rect 386 -1050 401 -1004
rect -280 -1116 -234 -1066
rect 325 -1067 401 -1050
rect 857 -1003 933 -990
rect 857 -1049 872 -1003
rect 918 -1049 933 -1003
rect 857 -1066 933 -1049
rect 340 -1116 386 -1067
rect -280 -1162 387 -1116
rect 865 -1233 925 -1066
rect -278 -1345 940 -1233
<< labels >>
flabel metal1 -165 -724 -116 -622 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 60 -725 109 -623 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 -282 -834 -231 -626 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 177 -832 228 -624 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 533 -947 747 -890 1 FreeSans 560 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 333 -1335 545 -1241 1 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional
flabel pwell -265 -1329 -118 -1244 1 FreeSans 368 0 0 0 VPW
port 7 nsew ground bidirectional
<< end >>
