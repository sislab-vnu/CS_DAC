magic
tech gf180mcuD
magscale 1 10
timestamp 1754896527
<< pwell >>
rect -356 -436 795 224
<< nmos >>
rect -200 -20 -144 24
rect -24 -20 32 24
rect 152 -20 208 24
rect 456 -20 512 24
rect 596 -20 652 24
rect -200 -248 -144 -160
rect -24 -248 336 -160
rect 596 -248 652 -160
<< ndiff >>
rect -124 24 -44 42
rect 52 25 132 42
rect 52 24 69 25
rect -246 -20 -200 24
rect -144 -20 -106 24
rect -124 -22 -106 -20
rect -60 -20 -24 24
rect 32 -20 69 24
rect -60 -22 -44 -20
rect -124 -38 -44 -22
rect 52 -21 69 -20
rect 115 24 132 25
rect 228 24 308 42
rect 115 -20 152 24
rect 208 -20 244 24
rect 115 -21 132 -20
rect 52 -38 132 -21
rect 228 -22 244 -20
rect 290 -22 308 24
rect 228 -38 308 -22
rect 364 25 436 38
rect 364 -21 377 25
rect 423 24 436 25
rect 423 -20 456 24
rect 512 -20 596 24
rect 652 -20 698 24
rect 423 -21 436 -20
rect 364 -34 436 -21
rect 532 -160 576 -20
rect -246 -248 -200 -160
rect -144 -186 -24 -160
rect -144 -232 -100 -186
rect -54 -232 -24 -186
rect -144 -248 -24 -232
rect 336 -248 596 -160
rect 652 -248 698 -160
<< ndiffc >>
rect -106 -22 -60 24
rect 69 -21 115 25
rect 244 -22 290 24
rect 377 -21 423 25
rect -100 -232 -54 -186
<< polysilicon >>
rect -36 147 44 164
rect -36 101 -19 147
rect 27 101 44 147
rect -36 84 44 101
rect 140 147 220 164
rect 140 101 157 147
rect 203 101 220 147
rect 140 84 220 101
rect 444 147 524 164
rect 444 101 461 147
rect 507 101 524 147
rect 444 84 524 101
rect -200 24 -144 70
rect -24 24 32 84
rect -200 -160 -144 -20
rect -24 -66 32 -20
rect 152 24 208 84
rect 152 -66 208 -20
rect 456 24 512 84
rect 596 24 652 70
rect 456 -104 512 -20
rect 300 -114 512 -104
rect -24 -140 512 -114
rect -24 -160 336 -140
rect 596 -160 652 -20
rect -200 -294 -144 -248
rect -24 -294 336 -248
rect 596 -294 652 -248
rect -212 -311 -132 -294
rect -212 -357 -195 -311
rect -149 -357 -132 -311
rect -212 -374 -132 -357
rect 584 -311 664 -294
rect 584 -357 601 -311
rect 647 -357 664 -311
rect 584 -374 664 -357
<< polycontact >>
rect -19 101 27 147
rect 157 101 203 147
rect 461 101 507 147
rect -195 -357 -149 -311
rect 601 -357 647 -311
<< metal1 >>
rect -34 147 42 162
rect -34 101 -19 147
rect 27 101 42 147
rect -34 86 42 101
rect 142 147 218 162
rect 142 101 157 147
rect 203 101 218 147
rect 142 86 218 101
rect 446 147 522 162
rect 446 101 461 147
rect 507 101 522 147
rect 446 86 522 101
rect -122 24 -46 40
rect -122 -22 -106 24
rect -60 -22 -46 24
rect -122 -36 -46 -22
rect 69 25 115 36
rect 69 -82 115 -21
rect 230 24 306 40
rect 230 -22 244 24
rect 290 -22 306 24
rect 230 -36 306 -22
rect 377 25 423 36
rect 377 -82 423 -21
rect 69 -128 423 -82
rect -114 -186 -38 -170
rect -114 -232 -100 -186
rect -54 -232 -38 -186
rect -114 -276 -38 -232
rect -266 -311 718 -276
rect -266 -357 -195 -311
rect -149 -357 601 -311
rect 647 -357 718 -311
rect -266 -396 718 -357
<< labels >>
flabel metal1 -34 86 42 162 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 142 86 218 162 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 -122 -36 -46 40 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 230 -36 306 40 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 446 86 522 162 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 -114 -396 -38 -232 1 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional
flabel pwell 479 -387 594 -286 1 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
<< end >>
