magic
tech gf180mcuD
magscale 1 10
timestamp 1755705775
<< pwell >>
rect -304 -185 1117 488
<< nmos >>
rect -166 240 -110 284
rect -14 240 42 284
rect 290 240 346 284
rect 466 240 522 284
rect 770 240 826 284
rect 928 240 984 284
rect -166 0 -110 90
rect 0 0 360 90
rect 452 0 812 90
rect 928 0 984 90
<< ndiff >>
rect 62 285 134 298
rect 62 284 75 285
rect -212 240 -166 284
rect -110 240 -14 284
rect 42 240 75 284
rect -80 90 -34 240
rect 62 239 75 240
rect 121 239 134 285
rect 62 226 134 239
rect 190 285 270 302
rect 190 239 207 285
rect 253 284 270 285
rect 366 287 446 304
rect 366 284 383 287
rect 253 240 290 284
rect 346 241 383 284
rect 429 284 446 287
rect 542 285 622 302
rect 542 284 559 285
rect 429 241 466 284
rect 346 240 466 241
rect 522 240 559 284
rect 253 239 270 240
rect 190 222 270 239
rect 366 224 446 240
rect 542 239 559 240
rect 605 239 622 285
rect 542 222 622 239
rect 678 285 750 298
rect 678 239 691 285
rect 737 284 750 285
rect 737 240 770 284
rect 826 240 928 284
rect 984 240 1030 284
rect 737 239 750 240
rect 678 226 750 239
rect 846 90 890 240
rect -212 0 -166 90
rect -110 0 0 90
rect 360 0 452 90
rect 812 0 928 90
rect 984 0 1030 90
rect 384 -56 428 0
rect 380 -66 432 -56
rect 366 -79 446 -66
rect 366 -125 381 -79
rect 427 -125 446 -79
rect 366 -138 446 -125
<< ndiffc >>
rect 75 239 121 285
rect 207 239 253 285
rect 383 241 429 287
rect 559 239 605 285
rect 691 239 737 285
rect 381 -125 427 -79
<< psubdiff >>
rect 679 -84 878 -71
rect 679 -130 753 -84
rect 799 -130 878 -84
rect 679 -143 878 -130
<< psubdiffcont >>
rect 753 -130 799 -84
<< polysilicon >>
rect -26 407 54 424
rect -26 361 -9 407
rect 37 361 54 407
rect -26 344 54 361
rect 278 407 358 424
rect 278 361 295 407
rect 341 361 358 407
rect 278 344 358 361
rect 454 407 534 424
rect 454 361 471 407
rect 517 361 534 407
rect 454 344 534 361
rect 758 407 838 424
rect 758 361 775 407
rect 821 361 838 407
rect 758 344 838 361
rect -166 284 -110 328
rect -14 284 42 344
rect -166 90 -110 240
rect -14 194 42 240
rect 290 284 346 344
rect 466 284 522 344
rect 290 194 346 240
rect 466 194 522 240
rect 770 284 826 344
rect 928 284 984 328
rect 770 194 826 240
rect 0 136 42 194
rect 324 136 488 146
rect 770 136 812 194
rect 0 110 812 136
rect 0 90 360 110
rect 452 90 812 110
rect 928 90 984 240
rect -166 -46 -110 0
rect 0 -46 360 0
rect -174 -59 -102 -46
rect 452 -46 812 0
rect 928 -46 984 0
rect -174 -105 -161 -59
rect -115 -105 -102 -59
rect 920 -59 992 -46
rect -174 -118 -102 -105
rect 920 -105 933 -59
rect 979 -105 992 -59
rect 920 -118 992 -105
<< polycontact >>
rect -9 361 37 407
rect 295 361 341 407
rect 471 361 517 407
rect 775 361 821 407
rect -161 -105 -115 -59
rect 933 -105 979 -59
<< metal1 >>
rect -24 407 52 422
rect -24 361 -9 407
rect 37 361 52 407
rect -24 346 52 361
rect 280 407 356 422
rect 280 361 295 407
rect 341 361 356 407
rect 280 346 356 361
rect 456 407 532 422
rect 456 361 471 407
rect 517 361 532 407
rect 456 346 532 361
rect 760 407 836 422
rect 760 361 775 407
rect 821 361 836 407
rect 760 346 836 361
rect 75 285 121 296
rect 75 168 121 239
rect 192 285 268 300
rect 192 239 207 285
rect 253 239 268 285
rect 192 224 268 239
rect 383 287 429 298
rect 383 168 429 241
rect 544 285 620 300
rect 544 239 559 285
rect 605 239 620 285
rect 544 224 620 239
rect 691 285 737 296
rect 691 168 737 239
rect 75 122 737 168
rect -200 -59 1016 -24
rect -200 -105 -161 -59
rect -115 -79 933 -59
rect -115 -105 381 -79
rect -200 -125 381 -105
rect 427 -84 933 -79
rect 427 -125 753 -84
rect -200 -130 753 -125
rect 799 -105 933 -84
rect 979 -105 1016 -59
rect 799 -130 1016 -105
rect -200 -144 1016 -130
<< labels >>
flabel metal1 280 346 356 422 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 456 346 532 422 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 192 224 268 300 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 544 224 620 300 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 760 346 836 422 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 -24 346 52 422 1 FreeSans 400 0 0 0 VBIAS
port 6 nsew power bidirectional
flabel metal1 -200 -144 1016 -24 1 FreeSans 400 0 0 0 VSS
port 7 n
<< end >>
