magic
tech gf180mcuD
magscale 1 10
timestamp 1756722462
<< nwell >>
rect 1344 67793 1400 67885
rect 6944 67793 7000 67885
rect 12544 67793 12600 67885
rect 18144 67793 18200 67885
rect 23744 67793 23800 67885
rect 29344 67793 29400 67885
rect 34944 67793 35000 67885
rect 1344 64209 1400 64301
rect 6944 64209 7000 64301
rect 12544 64209 12600 64301
rect 18144 64209 18200 64301
rect 23744 64209 23800 64301
rect 29344 64209 29400 64301
rect 34944 64209 35000 64301
rect 40544 64209 40600 64301
rect 1344 60625 1400 60717
rect 6944 60625 7000 60717
rect 12544 60625 12600 60717
rect 18144 60625 18200 60717
rect 23744 60625 23800 60717
rect 29344 60625 29400 60717
rect 34944 60625 35000 60717
rect 40544 60625 40600 60717
rect 1344 57041 1400 57133
rect 6944 57041 7000 57133
rect 12544 57041 12600 57133
rect 18144 57041 18200 57133
rect 23744 57041 23800 57133
rect 29344 57041 29400 57133
rect 34944 57041 35000 57133
rect 40544 57041 40600 57133
rect 1344 53457 1400 53549
rect 6944 53457 7000 53549
rect 12544 53457 12600 53549
rect 18144 53457 18200 53549
rect 23744 53457 23800 53549
rect 29344 53457 29400 53549
rect 34944 53457 35000 53549
rect 40544 53457 40600 53549
rect 1344 49873 1400 49965
rect 6944 49873 7000 49965
rect 12544 49873 12600 49965
rect 18144 49873 18200 49965
rect 23744 49873 23800 49965
rect 29344 49873 29400 49965
rect 34944 49873 35000 49965
rect 40544 49873 40600 49965
rect 1344 46289 1400 46381
rect 6944 46289 7000 46381
rect 12544 46289 12600 46381
rect 18144 46289 18200 46381
rect 23744 46289 23800 46381
rect 29344 46289 29400 46381
rect 34944 46289 35000 46381
rect 40544 46289 40600 46381
rect 1344 42705 1400 42737
rect 6944 42705 7000 42797
rect 12544 42705 12600 42797
rect 18144 42705 18200 42797
rect 23744 42705 23800 42797
rect 29344 42705 29400 42797
rect 34944 42705 35000 42797
<< metal1 >>
rect -952 70224 -784 70461
rect -952 70168 44240 70224
rect -952 70112 -112 70168
rect -56 70112 5488 70168
rect 5544 70112 11088 70168
rect 11144 70112 16688 70168
rect 16744 70112 22288 70168
rect 22344 70112 27888 70168
rect 27944 70112 33488 70168
rect 33544 70112 44240 70168
rect -952 70056 44240 70112
rect -952 66640 -784 70056
rect -168 69832 44240 69888
rect -168 69776 4467 69832
rect 4523 69776 10067 69832
rect 10123 69776 15667 69832
rect 15723 69776 21267 69832
rect 21323 69776 26867 69832
rect 26923 69776 32467 69832
rect 32523 69776 38067 69832
rect 38123 69776 44128 69832
rect 44184 69776 44240 69832
rect -168 69720 44240 69776
rect 44408 69552 44744 70565
rect -168 69384 44744 69552
rect -112 69259 -56 69272
rect -112 68834 -56 69203
rect 3985 69157 4041 69384
rect 4467 69256 4523 69272
rect 4467 69048 4523 69200
rect 5488 69259 5544 69272
rect 5488 68834 5544 69203
rect 9585 69157 9641 69384
rect 10067 69256 10123 69272
rect 10067 69048 10123 69200
rect 11088 69259 11144 69272
rect 11088 68834 11144 69203
rect 15185 69157 15241 69384
rect 15667 69256 15723 69272
rect 15667 69048 15723 69200
rect -112 68778 311 68834
rect 5488 68778 5911 68834
rect 11088 68778 11511 68834
rect 234 68234 290 68235
rect 238 68091 290 68234
rect 5838 68091 5890 68234
rect 11438 68091 11490 68247
rect 16520 67988 16576 69272
rect 16688 69259 16744 69272
rect 16688 68834 16744 69203
rect 20785 69157 20841 69384
rect 21267 69256 21323 69272
rect 21267 69048 21323 69200
rect 16688 68778 17111 68834
rect 17038 68091 17090 68247
rect 22120 67988 22176 69272
rect 22288 69259 22344 69272
rect 22288 68834 22344 69203
rect 26385 69157 26441 69384
rect 26867 69256 26923 69272
rect 26867 69048 26923 69200
rect 22288 68778 22711 68834
rect 22638 68091 22690 68247
rect 27720 67988 27776 69272
rect 27888 69259 27944 69272
rect 27888 68834 27944 69203
rect 31985 69157 32041 69384
rect 32467 69256 32523 69272
rect 32467 69048 32523 69200
rect 27888 68778 28311 68834
rect 28238 68091 28290 68247
rect 33320 67988 33376 69272
rect 33488 69259 33544 69272
rect 33488 68834 33544 69203
rect 37585 69157 37641 69384
rect 38067 69256 38123 69272
rect 38067 69048 38123 69200
rect 33488 68778 33911 68834
rect 33838 68091 33890 68247
rect 16520 67932 17092 67988
rect 22120 67932 22692 67988
rect 27720 67932 28292 67988
rect 33320 67932 33892 67988
rect -168 67312 44240 67368
rect -168 67256 4435 67312
rect 4491 67256 10035 67312
rect 10091 67256 15635 67312
rect 15691 67256 21235 67312
rect 21291 67256 26835 67312
rect 26891 67256 32435 67312
rect 32491 67256 38035 67312
rect 38091 67256 44128 67312
rect 44184 67256 44240 67312
rect -168 67200 44240 67256
rect -336 66976 44240 67032
rect -336 66920 -280 66976
rect -224 66920 1344 66976
rect 1400 66920 5320 66976
rect 5376 66920 6944 66976
rect 7000 66920 10920 66976
rect 10976 66920 12544 66976
rect 12600 66920 16520 66976
rect 16576 66920 18144 66976
rect 18200 66920 22120 66976
rect 22176 66920 23744 66976
rect 23800 66920 27720 66976
rect 27776 66920 29344 66976
rect 29400 66920 33320 66976
rect 33376 66920 34944 66976
rect 35000 66920 38920 66976
rect 38976 66920 44240 66976
rect -336 66864 44240 66920
rect -952 66584 44240 66640
rect -952 66528 -112 66584
rect -56 66528 5488 66584
rect 5544 66528 11088 66584
rect 11144 66528 16688 66584
rect 16744 66528 22288 66584
rect 22344 66528 27888 66584
rect 27944 66528 33488 66584
rect 33544 66528 39088 66584
rect 39144 66528 44240 66584
rect -952 66472 44240 66528
rect -952 63056 -784 66472
rect -168 66248 44240 66304
rect -168 66192 4467 66248
rect 4523 66192 10067 66248
rect 10123 66192 15667 66248
rect 15723 66192 21267 66248
rect 21323 66192 26867 66248
rect 26923 66192 32467 66248
rect 32523 66192 38067 66248
rect 38123 66192 43667 66248
rect 43723 66192 44128 66248
rect 44184 66192 44240 66248
rect -168 66136 44240 66192
rect 44408 65968 44744 69384
rect -168 65800 44744 65968
rect -280 65676 -224 65688
rect -280 64404 -224 65620
rect -112 65675 -56 65688
rect -112 65250 -56 65619
rect 3985 65573 4041 65800
rect 4467 65672 4523 65688
rect 4467 65464 4523 65616
rect 5320 65676 5376 65688
rect -112 65194 311 65250
rect 5320 64404 5376 65620
rect 5488 65675 5544 65688
rect 5488 65250 5544 65619
rect 9585 65573 9641 65800
rect 10067 65672 10123 65688
rect 10067 65464 10123 65616
rect 10920 65676 10976 65688
rect 5488 65194 5911 65250
rect 10920 64404 10976 65620
rect 11088 65675 11144 65688
rect 11088 65250 11144 65619
rect 15185 65573 15241 65800
rect 15667 65672 15723 65688
rect 15667 65464 15723 65616
rect 16520 65676 16576 65688
rect 11088 65194 11511 65250
rect 16520 64404 16576 65620
rect 16688 65675 16744 65688
rect 16688 65250 16744 65619
rect 20785 65573 20841 65800
rect 21267 65672 21323 65688
rect 21267 65464 21323 65616
rect 22120 65676 22176 65688
rect 16688 65194 17111 65250
rect 22120 64404 22176 65620
rect 22288 65675 22344 65688
rect 22288 65250 22344 65619
rect 26385 65573 26441 65800
rect 26867 65672 26923 65688
rect 26867 65464 26923 65616
rect 27720 65676 27776 65688
rect 22288 65194 22711 65250
rect 27720 64404 27776 65620
rect 27888 65675 27944 65688
rect 27888 65250 27944 65619
rect 31985 65573 32041 65800
rect 32467 65672 32523 65688
rect 32467 65464 32523 65616
rect 33320 65676 33376 65688
rect 27888 65194 28311 65250
rect 33320 64404 33376 65620
rect 33488 65675 33544 65688
rect 33488 65250 33544 65619
rect 37585 65573 37641 65800
rect 38067 65672 38123 65688
rect 38067 65464 38123 65616
rect 38920 65676 38976 65688
rect 33488 65194 33911 65250
rect 38920 64404 38976 65620
rect 39088 65675 39144 65688
rect 39088 65250 39144 65619
rect 43185 65573 43241 65800
rect 43667 65672 43723 65688
rect 43667 65464 43723 65616
rect 39088 65194 39511 65250
rect -280 64348 292 64404
rect 5320 64348 5892 64404
rect 10920 64348 11492 64404
rect 16520 64348 17092 64404
rect 22120 64348 22692 64404
rect 27720 64348 28292 64404
rect 33320 64348 33892 64404
rect 38920 64348 39492 64404
rect -168 63728 44240 63784
rect -168 63672 4435 63728
rect 4491 63672 10035 63728
rect 10091 63672 15635 63728
rect 15691 63672 21235 63728
rect 21291 63672 26835 63728
rect 26891 63672 32435 63728
rect 32491 63672 38035 63728
rect 38091 63672 43635 63728
rect 43691 63672 44128 63728
rect 44184 63672 44240 63728
rect -168 63616 44240 63672
rect -336 63392 44240 63448
rect -336 63336 -280 63392
rect -224 63336 1344 63392
rect 1400 63336 5320 63392
rect 5376 63336 6944 63392
rect 7000 63336 10920 63392
rect 10976 63336 12544 63392
rect 12600 63336 16520 63392
rect 16576 63336 18144 63392
rect 18200 63336 22120 63392
rect 22176 63336 23744 63392
rect 23800 63336 27720 63392
rect 27776 63336 29344 63392
rect 29400 63336 33320 63392
rect 33376 63336 34944 63392
rect 35000 63336 38920 63392
rect 38976 63336 40544 63392
rect 40600 63336 44240 63392
rect -336 63280 44240 63336
rect -952 63000 44240 63056
rect -952 62944 -112 63000
rect -56 62944 5488 63000
rect 5544 62944 11088 63000
rect 11144 62944 16688 63000
rect 16744 62944 22288 63000
rect 22344 62944 27888 63000
rect 27944 62944 33488 63000
rect 33544 62944 39088 63000
rect 39144 62944 44240 63000
rect -952 62888 44240 62944
rect -952 59472 -784 62888
rect -168 62664 44240 62720
rect -168 62608 4467 62664
rect 4523 62608 10067 62664
rect 10123 62608 15667 62664
rect 15723 62608 21267 62664
rect 21323 62608 26867 62664
rect 26923 62608 32467 62664
rect 32523 62608 38067 62664
rect 38123 62608 43667 62664
rect 43723 62608 44128 62664
rect 44184 62608 44240 62664
rect -168 62552 44240 62608
rect 44408 62384 44744 65800
rect -168 62216 44744 62384
rect -280 62092 -224 62104
rect -280 60820 -224 62036
rect -112 62091 -56 62104
rect -112 61666 -56 62035
rect 3985 61989 4041 62216
rect 4467 62088 4523 62104
rect 4467 61880 4523 62032
rect 5320 62092 5376 62104
rect -112 61610 311 61666
rect 5320 60820 5376 62036
rect 5488 62091 5544 62104
rect 5488 61666 5544 62035
rect 9585 61989 9641 62216
rect 10067 62088 10123 62104
rect 10067 61880 10123 62032
rect 10920 62092 10976 62104
rect 5488 61610 5911 61666
rect 10920 60820 10976 62036
rect 11088 62091 11144 62104
rect 11088 61666 11144 62035
rect 15185 61989 15241 62216
rect 15667 62088 15723 62104
rect 15667 61880 15723 62032
rect 16520 62092 16576 62104
rect 11088 61610 11511 61666
rect 16520 60820 16576 62036
rect 16688 62091 16744 62104
rect 16688 61666 16744 62035
rect 20785 61989 20841 62216
rect 21267 62088 21323 62104
rect 21267 61880 21323 62032
rect 22120 62092 22176 62104
rect 16688 61610 17111 61666
rect 22120 60820 22176 62036
rect 22288 62091 22344 62104
rect 22288 61666 22344 62035
rect 26385 61989 26441 62216
rect 26867 62088 26923 62104
rect 26867 61880 26923 62032
rect 27720 62092 27776 62104
rect 22288 61610 22711 61666
rect 27720 60820 27776 62036
rect 27888 62091 27944 62104
rect 27888 61666 27944 62035
rect 31985 61989 32041 62216
rect 32467 62088 32523 62104
rect 32467 61880 32523 62032
rect 33320 62092 33376 62104
rect 27888 61610 28311 61666
rect 33320 60820 33376 62036
rect 33488 62091 33544 62104
rect 33488 61666 33544 62035
rect 37585 61989 37641 62216
rect 38067 62088 38123 62104
rect 38067 61880 38123 62032
rect 38920 62092 38976 62104
rect 33488 61610 33911 61666
rect 38920 60820 38976 62036
rect 39088 62091 39144 62104
rect 39088 61666 39144 62035
rect 43185 61989 43241 62216
rect 43667 62088 43723 62104
rect 43667 61880 43723 62032
rect 39088 61610 39511 61666
rect -280 60764 292 60820
rect 5320 60764 5892 60820
rect 10920 60764 11492 60820
rect 16520 60764 17092 60820
rect 22120 60764 22692 60820
rect 27720 60764 28292 60820
rect 33320 60764 33892 60820
rect 38920 60764 39492 60820
rect -168 60144 44240 60200
rect -168 60088 4435 60144
rect 4491 60088 10035 60144
rect 10091 60088 15635 60144
rect 15691 60088 21235 60144
rect 21291 60088 26835 60144
rect 26891 60088 32435 60144
rect 32491 60088 38035 60144
rect 38091 60088 43635 60144
rect 43691 60088 44128 60144
rect 44184 60088 44240 60144
rect -168 60032 44240 60088
rect -336 59808 44240 59864
rect -336 59752 -280 59808
rect -224 59752 1344 59808
rect 1400 59752 5320 59808
rect 5376 59752 6944 59808
rect 7000 59752 10920 59808
rect 10976 59752 12544 59808
rect 12600 59752 16520 59808
rect 16576 59752 18144 59808
rect 18200 59752 22120 59808
rect 22176 59752 23744 59808
rect 23800 59752 27720 59808
rect 27776 59752 29344 59808
rect 29400 59752 33320 59808
rect 33376 59752 34944 59808
rect 35000 59752 38920 59808
rect 38976 59752 40544 59808
rect 40600 59752 44240 59808
rect -336 59696 44240 59752
rect -952 59416 44240 59472
rect -952 59360 -112 59416
rect -56 59360 5488 59416
rect 5544 59360 11088 59416
rect 11144 59360 16688 59416
rect 16744 59360 22288 59416
rect 22344 59360 27888 59416
rect 27944 59360 33488 59416
rect 33544 59360 39088 59416
rect 39144 59360 44240 59416
rect -952 59304 44240 59360
rect -952 55888 -784 59304
rect -168 59080 44240 59136
rect -168 59024 4467 59080
rect 4523 59024 10067 59080
rect 10123 59024 15667 59080
rect 15723 59024 21267 59080
rect 21323 59024 26867 59080
rect 26923 59024 32467 59080
rect 32523 59024 38067 59080
rect 38123 59024 43667 59080
rect 43723 59024 44128 59080
rect 44184 59024 44240 59080
rect -168 58968 44240 59024
rect 44408 58800 44744 62216
rect -168 58632 44744 58800
rect -280 58508 -224 58520
rect -280 57236 -224 58452
rect -112 58507 -56 58520
rect -112 58082 -56 58451
rect 3985 58405 4041 58632
rect 4467 58504 4523 58520
rect 4467 58296 4523 58448
rect 5320 58508 5376 58520
rect -112 58026 311 58082
rect 5320 57236 5376 58452
rect 5488 58507 5544 58520
rect 5488 58082 5544 58451
rect 9585 58405 9641 58632
rect 10067 58504 10123 58520
rect 10067 58296 10123 58448
rect 10920 58508 10976 58520
rect 5488 58026 5911 58082
rect 10920 57236 10976 58452
rect 11088 58507 11144 58520
rect 11088 58082 11144 58451
rect 15185 58405 15241 58632
rect 15667 58504 15723 58520
rect 15667 58296 15723 58448
rect 16520 58508 16576 58520
rect 11088 58026 11511 58082
rect 16520 57236 16576 58452
rect 16688 58507 16744 58520
rect 16688 58082 16744 58451
rect 20785 58405 20841 58632
rect 21267 58504 21323 58520
rect 21267 58296 21323 58448
rect 22120 58508 22176 58520
rect 16688 58026 17111 58082
rect 22120 57236 22176 58452
rect 22288 58507 22344 58520
rect 22288 58082 22344 58451
rect 26385 58405 26441 58632
rect 26867 58504 26923 58520
rect 26867 58296 26923 58448
rect 27720 58508 27776 58520
rect 22288 58026 22711 58082
rect 27720 57236 27776 58452
rect 27888 58507 27944 58520
rect 27888 58082 27944 58451
rect 31985 58405 32041 58632
rect 32467 58504 32523 58520
rect 32467 58296 32523 58448
rect 33320 58508 33376 58520
rect 27888 58026 28311 58082
rect 33320 57236 33376 58452
rect 33488 58507 33544 58520
rect 33488 58082 33544 58451
rect 37585 58405 37641 58632
rect 38067 58504 38123 58520
rect 38067 58296 38123 58448
rect 38920 58508 38976 58520
rect 33488 58026 33911 58082
rect 38920 57236 38976 58452
rect 39088 58507 39144 58520
rect 39088 58082 39144 58451
rect 43185 58405 43241 58632
rect 43667 58504 43723 58520
rect 43667 58296 43723 58448
rect 39088 58026 39511 58082
rect -280 57180 292 57236
rect 5320 57180 5892 57236
rect 10920 57180 11492 57236
rect 16520 57180 17092 57236
rect 22120 57180 22692 57236
rect 27720 57180 28292 57236
rect 33320 57180 33892 57236
rect 38920 57180 39492 57236
rect -168 56560 44240 56616
rect -168 56504 4435 56560
rect 4491 56504 10035 56560
rect 10091 56504 15635 56560
rect 15691 56504 21235 56560
rect 21291 56504 26835 56560
rect 26891 56504 32435 56560
rect 32491 56504 38035 56560
rect 38091 56504 43635 56560
rect 43691 56504 44128 56560
rect 44184 56504 44240 56560
rect -168 56448 44240 56504
rect -336 56224 44240 56280
rect -336 56168 -280 56224
rect -224 56168 1344 56224
rect 1400 56168 5320 56224
rect 5376 56168 6944 56224
rect 7000 56168 10920 56224
rect 10976 56168 12544 56224
rect 12600 56168 16520 56224
rect 16576 56168 18144 56224
rect 18200 56168 22120 56224
rect 22176 56168 23744 56224
rect 23800 56168 27720 56224
rect 27776 56168 29344 56224
rect 29400 56168 33320 56224
rect 33376 56168 34944 56224
rect 35000 56168 38920 56224
rect 38976 56168 40544 56224
rect 40600 56168 44240 56224
rect -336 56112 44240 56168
rect -952 55832 44240 55888
rect -952 55776 -112 55832
rect -56 55776 5488 55832
rect 5544 55776 11088 55832
rect 11144 55776 16688 55832
rect 16744 55776 22288 55832
rect 22344 55776 27888 55832
rect 27944 55776 33488 55832
rect 33544 55776 39088 55832
rect 39144 55776 44240 55832
rect -952 55720 44240 55776
rect -952 52304 -784 55720
rect -168 55496 44240 55552
rect -168 55440 4467 55496
rect 4523 55440 10067 55496
rect 10123 55440 15667 55496
rect 15723 55440 21267 55496
rect 21323 55440 26867 55496
rect 26923 55440 32467 55496
rect 32523 55440 38067 55496
rect 38123 55440 43667 55496
rect 43723 55440 44128 55496
rect 44184 55440 44240 55496
rect -168 55384 44240 55440
rect 44408 55216 44744 58632
rect -168 55048 44744 55216
rect -280 54924 -224 54936
rect -280 53652 -224 54868
rect -112 54923 -56 54936
rect -112 54498 -56 54867
rect 3985 54821 4041 55048
rect 4467 54920 4523 54936
rect 4467 54712 4523 54864
rect 5320 54924 5376 54936
rect -112 54442 311 54498
rect 5320 53652 5376 54868
rect 5488 54923 5544 54936
rect 5488 54498 5544 54867
rect 9585 54821 9641 55048
rect 10067 54920 10123 54936
rect 10067 54712 10123 54864
rect 10920 54924 10976 54936
rect 5488 54442 5911 54498
rect 10920 53652 10976 54868
rect 11088 54923 11144 54936
rect 11088 54498 11144 54867
rect 15185 54821 15241 55048
rect 15667 54920 15723 54936
rect 15667 54712 15723 54864
rect 16520 54924 16576 54936
rect 11088 54442 11511 54498
rect 16520 53652 16576 54868
rect 16688 54923 16744 54936
rect 16688 54498 16744 54867
rect 20785 54821 20841 55048
rect 21267 54920 21323 54936
rect 21267 54712 21323 54864
rect 22120 54924 22176 54936
rect 16688 54442 17111 54498
rect 22120 53652 22176 54868
rect 22288 54923 22344 54936
rect 22288 54498 22344 54867
rect 26385 54821 26441 55048
rect 26867 54920 26923 54936
rect 26867 54712 26923 54864
rect 27720 54924 27776 54936
rect 22288 54442 22711 54498
rect 27720 53652 27776 54868
rect 27888 54923 27944 54936
rect 27888 54498 27944 54867
rect 31985 54821 32041 55048
rect 32467 54920 32523 54936
rect 32467 54712 32523 54864
rect 33320 54924 33376 54936
rect 27888 54442 28311 54498
rect 33320 53652 33376 54868
rect 33488 54923 33544 54936
rect 33488 54498 33544 54867
rect 37585 54821 37641 55048
rect 38067 54920 38123 54936
rect 38067 54712 38123 54864
rect 38920 54924 38976 54936
rect 33488 54442 33911 54498
rect 38920 53652 38976 54868
rect 39088 54923 39144 54936
rect 39088 54498 39144 54867
rect 43185 54821 43241 55048
rect 43667 54920 43723 54936
rect 43667 54712 43723 54864
rect 39088 54442 39511 54498
rect -280 53596 292 53652
rect 5320 53596 5892 53652
rect 10920 53596 11492 53652
rect 16520 53596 17092 53652
rect 22120 53596 22692 53652
rect 27720 53596 28292 53652
rect 33320 53596 33892 53652
rect 38920 53596 39492 53652
rect -168 52976 44240 53032
rect -168 52920 4435 52976
rect 4491 52920 10035 52976
rect 10091 52920 15635 52976
rect 15691 52920 21235 52976
rect 21291 52920 26835 52976
rect 26891 52920 32435 52976
rect 32491 52920 38035 52976
rect 38091 52920 43635 52976
rect 43691 52920 44128 52976
rect 44184 52920 44240 52976
rect -168 52864 44240 52920
rect -336 52640 44240 52696
rect -336 52584 -280 52640
rect -224 52584 1344 52640
rect 1400 52584 5320 52640
rect 5376 52584 6944 52640
rect 7000 52584 10920 52640
rect 10976 52584 12544 52640
rect 12600 52584 16520 52640
rect 16576 52584 18144 52640
rect 18200 52584 22120 52640
rect 22176 52584 23744 52640
rect 23800 52584 27720 52640
rect 27776 52584 29344 52640
rect 29400 52584 33320 52640
rect 33376 52584 34944 52640
rect 35000 52584 38920 52640
rect 38976 52584 40544 52640
rect 40600 52584 44240 52640
rect -336 52528 44240 52584
rect -952 52248 44240 52304
rect -952 52192 -112 52248
rect -56 52192 5488 52248
rect 5544 52192 11088 52248
rect 11144 52192 16688 52248
rect 16744 52192 22288 52248
rect 22344 52192 27888 52248
rect 27944 52192 33488 52248
rect 33544 52192 39088 52248
rect 39144 52192 44240 52248
rect -952 52136 44240 52192
rect -952 48720 -784 52136
rect -168 51912 44240 51968
rect -168 51856 4467 51912
rect 4523 51856 10067 51912
rect 10123 51856 15667 51912
rect 15723 51856 21267 51912
rect 21323 51856 26867 51912
rect 26923 51856 32467 51912
rect 32523 51856 38067 51912
rect 38123 51856 43667 51912
rect 43723 51856 44128 51912
rect 44184 51856 44240 51912
rect -168 51800 44240 51856
rect 44408 51632 44744 55048
rect -168 51464 44744 51632
rect -280 51340 -224 51352
rect -280 50068 -224 51284
rect -112 51339 -56 51352
rect -112 50914 -56 51283
rect 3985 51237 4041 51464
rect 4467 51336 4523 51352
rect 4467 51128 4523 51280
rect 5320 51340 5376 51352
rect -112 50858 311 50914
rect 5320 50068 5376 51284
rect 5488 51339 5544 51352
rect 5488 50914 5544 51283
rect 9585 51237 9641 51464
rect 10067 51336 10123 51352
rect 10067 51128 10123 51280
rect 10920 51340 10976 51352
rect 5488 50858 5911 50914
rect 10920 50068 10976 51284
rect 11088 51339 11144 51352
rect 11088 50914 11144 51283
rect 15185 51237 15241 51464
rect 15667 51336 15723 51352
rect 15667 51128 15723 51280
rect 16520 51340 16576 51352
rect 11088 50858 11511 50914
rect 16520 50068 16576 51284
rect 16688 51339 16744 51352
rect 16688 50914 16744 51283
rect 20785 51237 20841 51464
rect 21267 51336 21323 51352
rect 21267 51128 21323 51280
rect 22120 51340 22176 51352
rect 16688 50858 17111 50914
rect 22120 50068 22176 51284
rect 22288 51339 22344 51352
rect 22288 50914 22344 51283
rect 26385 51237 26441 51464
rect 26867 51336 26923 51352
rect 26867 51128 26923 51280
rect 27720 51340 27776 51352
rect 22288 50858 22711 50914
rect 27720 50068 27776 51284
rect 27888 51339 27944 51352
rect 27888 50914 27944 51283
rect 31985 51237 32041 51464
rect 32467 51336 32523 51352
rect 32467 51128 32523 51280
rect 33320 51340 33376 51352
rect 27888 50858 28311 50914
rect 33320 50068 33376 51284
rect 33488 51339 33544 51352
rect 33488 50914 33544 51283
rect 37585 51237 37641 51464
rect 38067 51336 38123 51352
rect 38067 51128 38123 51280
rect 38920 51340 38976 51352
rect 33488 50858 33911 50914
rect 38920 50068 38976 51284
rect 39088 51339 39144 51352
rect 39088 50914 39144 51283
rect 43185 51237 43241 51464
rect 43667 51336 43723 51352
rect 43667 51128 43723 51280
rect 39088 50858 39511 50914
rect -280 50012 292 50068
rect 5320 50012 5892 50068
rect 10920 50012 11492 50068
rect 16520 50012 17092 50068
rect 22120 50012 22692 50068
rect 27720 50012 28292 50068
rect 33320 50012 33892 50068
rect 38920 50012 39492 50068
rect -168 49392 44240 49448
rect -168 49336 4435 49392
rect 4491 49336 10035 49392
rect 10091 49336 15635 49392
rect 15691 49336 21235 49392
rect 21291 49336 26835 49392
rect 26891 49336 32435 49392
rect 32491 49336 38035 49392
rect 38091 49336 43635 49392
rect 43691 49336 44128 49392
rect 44184 49336 44240 49392
rect -168 49280 44240 49336
rect -336 49056 44240 49112
rect -336 49000 -280 49056
rect -224 49000 1344 49056
rect 1400 49000 5320 49056
rect 5376 49000 6944 49056
rect 7000 49000 10920 49056
rect 10976 49000 12544 49056
rect 12600 49000 16520 49056
rect 16576 49000 18144 49056
rect 18200 49000 22120 49056
rect 22176 49000 23744 49056
rect 23800 49000 27720 49056
rect 27776 49000 29344 49056
rect 29400 49000 33320 49056
rect 33376 49000 34944 49056
rect 35000 49000 38920 49056
rect 38976 49000 40544 49056
rect 40600 49000 44240 49056
rect -336 48944 44240 49000
rect -952 48664 44240 48720
rect -952 48608 -112 48664
rect -56 48608 5488 48664
rect 5544 48608 11088 48664
rect 11144 48608 16688 48664
rect 16744 48608 22288 48664
rect 22344 48608 27888 48664
rect 27944 48608 33488 48664
rect 33544 48608 39088 48664
rect 39144 48608 44240 48664
rect -952 48552 44240 48608
rect -952 45136 -784 48552
rect -168 48328 44240 48384
rect -168 48272 4467 48328
rect 4523 48272 10067 48328
rect 10123 48272 15667 48328
rect 15723 48272 21267 48328
rect 21323 48272 26867 48328
rect 26923 48272 32467 48328
rect 32523 48272 38067 48328
rect 38123 48272 43667 48328
rect 43723 48272 44128 48328
rect 44184 48272 44240 48328
rect -168 48216 44240 48272
rect 44408 48048 44744 51464
rect -168 47880 44744 48048
rect -280 47755 -224 47768
rect -280 46484 -224 47699
rect -112 47755 -56 47768
rect -112 47330 -56 47699
rect 3985 47653 4041 47880
rect 4467 47752 4523 47768
rect 4467 47544 4523 47696
rect 5320 47756 5376 47768
rect -112 47274 311 47330
rect 5320 46484 5376 47700
rect 5488 47755 5544 47768
rect 5488 47330 5544 47699
rect 9585 47653 9641 47880
rect 10067 47752 10123 47768
rect 10067 47544 10123 47696
rect 10920 47756 10976 47768
rect 5488 47274 5911 47330
rect 10920 46484 10976 47700
rect 11088 47755 11144 47768
rect 11088 47330 11144 47699
rect 15185 47653 15241 47880
rect 15667 47752 15723 47768
rect 15667 47544 15723 47696
rect 16520 47755 16576 47768
rect 11088 47274 11511 47330
rect 16520 46484 16576 47699
rect 16688 47755 16744 47768
rect 16688 47330 16744 47699
rect 20785 47653 20841 47880
rect 21267 47752 21323 47768
rect 21267 47544 21323 47696
rect 22120 47756 22176 47768
rect 16688 47274 17111 47330
rect 22120 46484 22176 47700
rect 22288 47755 22344 47768
rect 22288 47330 22344 47699
rect 26385 47653 26441 47880
rect 26867 47752 26923 47768
rect 26867 47544 26923 47696
rect 27720 47756 27776 47768
rect 22288 47274 22711 47330
rect 27720 46484 27776 47700
rect 27888 47755 27944 47768
rect 27888 47330 27944 47699
rect 31985 47653 32041 47880
rect 32467 47752 32523 47768
rect 32467 47544 32523 47696
rect 33320 47756 33376 47768
rect 27888 47274 28311 47330
rect 33320 46484 33376 47700
rect 33488 47755 33544 47768
rect 33488 47330 33544 47699
rect 37585 47653 37641 47880
rect 38067 47752 38123 47768
rect 38067 47544 38123 47696
rect 38920 47756 38976 47768
rect 33488 47274 33911 47330
rect 38920 46484 38976 47700
rect 39088 47755 39144 47768
rect 39088 47330 39144 47699
rect 43185 47653 43241 47880
rect 43667 47752 43723 47768
rect 43667 47544 43723 47696
rect 39088 47274 39511 47330
rect -280 46428 292 46484
rect 5320 46428 5892 46484
rect 10920 46428 11492 46484
rect 16520 46428 17092 46484
rect 22120 46428 22692 46484
rect 27720 46428 28292 46484
rect 33320 46428 33892 46484
rect 38920 46428 39492 46484
rect -168 45808 44240 45864
rect -168 45752 4435 45808
rect 4491 45752 10035 45808
rect 10091 45752 15635 45808
rect 15691 45752 21235 45808
rect 21291 45752 26835 45808
rect 26891 45752 32435 45808
rect 32491 45752 38035 45808
rect 38091 45752 43635 45808
rect 43691 45752 44128 45808
rect 44184 45752 44240 45808
rect -168 45696 44240 45752
rect -336 45472 44240 45528
rect -336 45416 -280 45472
rect -224 45416 1344 45472
rect 1400 45416 5320 45472
rect 5376 45416 6944 45472
rect 7000 45416 10920 45472
rect 10976 45416 12544 45472
rect 12600 45416 16520 45472
rect 16576 45416 18144 45472
rect 18200 45416 22120 45472
rect 22176 45416 23744 45472
rect 23800 45416 27720 45472
rect 27776 45416 29344 45472
rect 29400 45416 33320 45472
rect 33376 45416 34944 45472
rect 35000 45416 38920 45472
rect 38976 45416 40544 45472
rect 40600 45416 44240 45472
rect -336 45360 44240 45416
rect -952 45080 44240 45136
rect -952 45024 -112 45080
rect -56 45024 5488 45080
rect 5544 45024 11088 45080
rect 11144 45024 16688 45080
rect 16744 45024 22288 45080
rect 22344 45024 27888 45080
rect 27944 45024 33488 45080
rect 33544 45024 39088 45080
rect 39144 45024 44240 45080
rect -952 44968 44240 45024
rect -952 41776 -784 44968
rect -168 44744 44240 44800
rect -168 44688 4467 44744
rect 4523 44688 10067 44744
rect 10123 44688 15667 44744
rect 15723 44688 21267 44744
rect 21323 44688 26867 44744
rect 26923 44688 32467 44744
rect 32523 44688 38067 44744
rect 38123 44688 43667 44744
rect 43723 44688 44128 44744
rect 44184 44688 44240 44744
rect -168 44632 44240 44688
rect 44408 44464 44744 47880
rect -168 44296 44744 44464
rect -280 44172 -224 44184
rect -280 42896 -224 44116
rect -112 44171 -56 44184
rect -112 43746 -56 44115
rect 3985 44069 4041 44296
rect 4467 44168 4523 44184
rect 4467 43960 4523 44112
rect 5320 44172 5376 44184
rect -112 43690 311 43746
rect 5320 42896 5376 44116
rect 5488 44171 5544 44184
rect 5488 43746 5544 44115
rect 9585 44069 9641 44296
rect 10067 44168 10123 44184
rect 10067 43960 10123 44112
rect 10920 44172 10976 44184
rect 5488 43690 5911 43746
rect 10920 42896 10976 44116
rect 11088 44171 11144 44184
rect 11088 43746 11144 44115
rect 15185 44069 15241 44296
rect 15667 44168 15723 44184
rect 15667 43960 15723 44112
rect 16520 44172 16576 44184
rect 11088 43690 11511 43746
rect 16520 42896 16576 44116
rect 16688 44171 16744 44184
rect 16688 43746 16744 44115
rect 20785 44069 20841 44296
rect 21267 44168 21323 44184
rect 21267 43960 21323 44112
rect 22120 44172 22176 44184
rect 16688 43690 17111 43746
rect 22120 42896 22176 44116
rect 22288 44171 22344 44184
rect 22288 43746 22344 44115
rect 26385 44069 26441 44296
rect 26867 44168 26923 44184
rect 26867 43960 26923 44112
rect 27720 44172 27776 44184
rect 22288 43690 22711 43746
rect 27720 42896 27776 44116
rect 27888 44171 27944 44184
rect 27888 43746 27944 44115
rect 31985 44069 32041 44296
rect 32467 44168 32523 44184
rect 32467 43960 32523 44112
rect 33320 44172 33376 44184
rect 27888 43690 28311 43746
rect 33320 42896 33376 44116
rect 33488 44171 33544 44184
rect 33488 43746 33544 44115
rect 37585 44069 37641 44296
rect 38067 44168 38123 44184
rect 38067 43960 38123 44112
rect 38920 44172 38976 44184
rect 33488 43690 33911 43746
rect 38920 42896 38976 44116
rect 39088 44171 39144 44184
rect 39088 43746 39144 44115
rect 43185 44051 43241 44296
rect 43667 44172 43723 44184
rect 43667 44008 43723 44116
rect 39088 43690 39604 43746
rect -280 42840 280 42896
rect 5320 42840 5890 42896
rect 10920 42840 11463 42896
rect 16520 42840 17079 42896
rect 22120 42840 22690 42896
rect 27720 42840 28261 42896
rect 33320 42839 33839 42896
rect 38920 42840 39446 42896
rect -168 42224 44240 42280
rect -168 42168 4435 42224
rect 4491 42168 10035 42224
rect 10091 42168 15635 42224
rect 15691 42168 21235 42224
rect 21291 42168 26835 42224
rect 26891 42168 32435 42224
rect 32491 42168 38035 42224
rect 38091 42168 43635 42224
rect 43691 42168 44128 42224
rect 44184 42168 44240 42224
rect -168 42112 44240 42168
rect 44408 41776 44744 44296
rect 44912 69832 45248 70565
rect 44912 69776 45024 69832
rect 45136 69776 45248 69832
rect 44912 66248 45248 69776
rect 44912 66192 45024 66248
rect 45136 66192 45248 66248
rect 44912 62664 45248 66192
rect 44912 62608 45024 62664
rect 45136 62608 45248 62664
rect 44912 59080 45248 62608
rect 44912 59024 45024 59080
rect 45136 59024 45248 59080
rect 44912 55496 45248 59024
rect 44912 55440 45024 55496
rect 45136 55440 45248 55496
rect 44912 51912 45248 55440
rect 44912 51856 45024 51912
rect 45136 51856 45248 51912
rect 44912 48328 45248 51856
rect 44912 48272 45024 48328
rect 45136 48272 45248 48328
rect 44912 44744 45248 48272
rect 44912 44688 45024 44744
rect 45136 44688 45248 44744
rect 44912 41776 45248 44688
rect 45416 67312 45752 70565
rect 45416 67256 45499 67312
rect 45611 67256 45752 67312
rect 45416 63728 45752 67256
rect 45416 63672 45497 63728
rect 45609 63672 45752 63728
rect 45416 60144 45752 63672
rect 45416 60088 45499 60144
rect 45611 60088 45752 60144
rect 45416 56560 45752 60088
rect 45416 56504 45497 56560
rect 45609 56504 45752 56560
rect 45416 52976 45752 56504
rect 45416 52920 45498 52976
rect 45610 52920 45752 52976
rect 45416 49392 45752 52920
rect 45416 49336 45500 49392
rect 45612 49336 45752 49392
rect 45416 45808 45752 49336
rect 45416 45752 45497 45808
rect 45609 45752 45752 45808
rect 45416 42224 45752 45752
rect 45416 42168 45498 42224
rect 45610 42168 45752 42224
rect 45416 41776 45752 42168
<< via1 >>
rect -112 70112 -56 70168
rect 5488 70112 5544 70168
rect 11088 70112 11144 70168
rect 16688 70112 16744 70168
rect 22288 70112 22344 70168
rect 27888 70112 27944 70168
rect 33488 70112 33544 70168
rect 4467 69776 4523 69832
rect 10067 69776 10123 69832
rect 15667 69776 15723 69832
rect 21267 69776 21323 69832
rect 26867 69776 26923 69832
rect 32467 69776 32523 69832
rect 38067 69776 38123 69832
rect 44128 69776 44184 69832
rect -112 69203 -56 69259
rect 4467 69200 4523 69256
rect 5488 69203 5544 69259
rect 10067 69200 10123 69256
rect 11088 69203 11144 69259
rect 15667 69200 15723 69256
rect 16688 69203 16744 69259
rect 21267 69200 21323 69256
rect 22288 69203 22344 69259
rect 26867 69200 26923 69256
rect 27888 69203 27944 69259
rect 32467 69200 32523 69256
rect 33488 69203 33544 69259
rect 38067 69200 38123 69256
rect 1667 67874 1723 67930
rect 7267 67874 7323 67930
rect 12867 67874 12923 67930
rect 18467 67874 18523 67930
rect 24067 67874 24123 67930
rect 29667 67874 29723 67930
rect 35267 67874 35323 67930
rect 448 67648 504 67704
rect 6048 67648 6104 67704
rect 11648 67648 11704 67704
rect 17248 67648 17304 67704
rect 22848 67648 22904 67704
rect 28448 67648 28504 67704
rect 34048 67648 34104 67704
rect 4435 67256 4491 67312
rect 10035 67256 10091 67312
rect 15635 67256 15691 67312
rect 21235 67256 21291 67312
rect 26835 67256 26891 67312
rect 32435 67256 32491 67312
rect 38035 67256 38091 67312
rect 44128 67256 44184 67312
rect -280 66920 -224 66976
rect 1344 66920 1400 66976
rect 5320 66920 5376 66976
rect 6944 66920 7000 66976
rect 10920 66920 10976 66976
rect 12544 66920 12600 66976
rect 16520 66920 16576 66976
rect 18144 66920 18200 66976
rect 22120 66920 22176 66976
rect 23744 66920 23800 66976
rect 27720 66920 27776 66976
rect 29344 66920 29400 66976
rect 33320 66920 33376 66976
rect 34944 66920 35000 66976
rect 38920 66920 38976 66976
rect -112 66528 -56 66584
rect 5488 66528 5544 66584
rect 11088 66528 11144 66584
rect 16688 66528 16744 66584
rect 22288 66528 22344 66584
rect 27888 66528 27944 66584
rect 33488 66528 33544 66584
rect 39088 66528 39144 66584
rect 4467 66192 4523 66248
rect 10067 66192 10123 66248
rect 15667 66192 15723 66248
rect 21267 66192 21323 66248
rect 26867 66192 26923 66248
rect 32467 66192 32523 66248
rect 38067 66192 38123 66248
rect 43667 66192 43723 66248
rect 44128 66192 44184 66248
rect -280 65620 -224 65676
rect -112 65619 -56 65675
rect 4467 65616 4523 65672
rect 5320 65620 5376 65676
rect 5488 65619 5544 65675
rect 10067 65616 10123 65672
rect 10920 65620 10976 65676
rect 11088 65619 11144 65675
rect 15667 65616 15723 65672
rect 16520 65620 16576 65676
rect 16688 65619 16744 65675
rect 21267 65616 21323 65672
rect 22120 65620 22176 65676
rect 22288 65619 22344 65675
rect 26867 65616 26923 65672
rect 27720 65620 27776 65676
rect 27888 65619 27944 65675
rect 32467 65616 32523 65672
rect 33320 65620 33376 65676
rect 33488 65619 33544 65675
rect 38067 65616 38123 65672
rect 38920 65620 38976 65676
rect 39088 65619 39144 65675
rect 43667 65616 43723 65672
rect 1667 64290 1723 64346
rect 7267 64290 7323 64346
rect 12867 64290 12923 64346
rect 18467 64290 18523 64346
rect 24067 64290 24123 64346
rect 29667 64290 29723 64346
rect 35267 64290 35323 64346
rect 40867 64290 40923 64346
rect 448 64064 504 64120
rect 6048 64064 6104 64120
rect 11648 64064 11704 64120
rect 17248 64064 17304 64120
rect 22848 64064 22904 64120
rect 28448 64064 28504 64120
rect 34048 64064 34104 64120
rect 39648 64064 39704 64120
rect 4435 63672 4491 63728
rect 10035 63672 10091 63728
rect 15635 63672 15691 63728
rect 21235 63672 21291 63728
rect 26835 63672 26891 63728
rect 32435 63672 32491 63728
rect 38035 63672 38091 63728
rect 43635 63672 43691 63728
rect 44128 63672 44184 63728
rect -280 63336 -224 63392
rect 1344 63336 1400 63392
rect 5320 63336 5376 63392
rect 6944 63336 7000 63392
rect 10920 63336 10976 63392
rect 12544 63336 12600 63392
rect 16520 63336 16576 63392
rect 18144 63336 18200 63392
rect 22120 63336 22176 63392
rect 23744 63336 23800 63392
rect 27720 63336 27776 63392
rect 29344 63336 29400 63392
rect 33320 63336 33376 63392
rect 34944 63336 35000 63392
rect 38920 63336 38976 63392
rect 40544 63336 40600 63392
rect -112 62944 -56 63000
rect 5488 62944 5544 63000
rect 11088 62944 11144 63000
rect 16688 62944 16744 63000
rect 22288 62944 22344 63000
rect 27888 62944 27944 63000
rect 33488 62944 33544 63000
rect 39088 62944 39144 63000
rect 4467 62608 4523 62664
rect 10067 62608 10123 62664
rect 15667 62608 15723 62664
rect 21267 62608 21323 62664
rect 26867 62608 26923 62664
rect 32467 62608 32523 62664
rect 38067 62608 38123 62664
rect 43667 62608 43723 62664
rect 44128 62608 44184 62664
rect -280 62036 -224 62092
rect -112 62035 -56 62091
rect 4467 62032 4523 62088
rect 5320 62036 5376 62092
rect 5488 62035 5544 62091
rect 10067 62032 10123 62088
rect 10920 62036 10976 62092
rect 11088 62035 11144 62091
rect 15667 62032 15723 62088
rect 16520 62036 16576 62092
rect 16688 62035 16744 62091
rect 21267 62032 21323 62088
rect 22120 62036 22176 62092
rect 22288 62035 22344 62091
rect 26867 62032 26923 62088
rect 27720 62036 27776 62092
rect 27888 62035 27944 62091
rect 32467 62032 32523 62088
rect 33320 62036 33376 62092
rect 33488 62035 33544 62091
rect 38067 62032 38123 62088
rect 38920 62036 38976 62092
rect 39088 62035 39144 62091
rect 43667 62032 43723 62088
rect 1667 60706 1723 60762
rect 7267 60706 7323 60762
rect 12867 60706 12923 60762
rect 18467 60706 18523 60762
rect 24067 60706 24123 60762
rect 29667 60706 29723 60762
rect 35267 60706 35323 60762
rect 40867 60706 40923 60762
rect 448 60480 504 60536
rect 6048 60480 6104 60536
rect 11648 60480 11704 60536
rect 17248 60480 17304 60536
rect 22848 60480 22904 60536
rect 28448 60480 28504 60536
rect 34048 60480 34104 60536
rect 39648 60480 39704 60536
rect 4435 60088 4491 60144
rect 10035 60088 10091 60144
rect 15635 60088 15691 60144
rect 21235 60088 21291 60144
rect 26835 60088 26891 60144
rect 32435 60088 32491 60144
rect 38035 60088 38091 60144
rect 43635 60088 43691 60144
rect 44128 60088 44184 60144
rect -280 59752 -224 59808
rect 1344 59752 1400 59808
rect 5320 59752 5376 59808
rect 6944 59752 7000 59808
rect 10920 59752 10976 59808
rect 12544 59752 12600 59808
rect 16520 59752 16576 59808
rect 18144 59752 18200 59808
rect 22120 59752 22176 59808
rect 23744 59752 23800 59808
rect 27720 59752 27776 59808
rect 29344 59752 29400 59808
rect 33320 59752 33376 59808
rect 34944 59752 35000 59808
rect 38920 59752 38976 59808
rect 40544 59752 40600 59808
rect -112 59360 -56 59416
rect 5488 59360 5544 59416
rect 11088 59360 11144 59416
rect 16688 59360 16744 59416
rect 22288 59360 22344 59416
rect 27888 59360 27944 59416
rect 33488 59360 33544 59416
rect 39088 59360 39144 59416
rect 4467 59024 4523 59080
rect 10067 59024 10123 59080
rect 15667 59024 15723 59080
rect 21267 59024 21323 59080
rect 26867 59024 26923 59080
rect 32467 59024 32523 59080
rect 38067 59024 38123 59080
rect 43667 59024 43723 59080
rect 44128 59024 44184 59080
rect -280 58452 -224 58508
rect -112 58451 -56 58507
rect 4467 58448 4523 58504
rect 5320 58452 5376 58508
rect 5488 58451 5544 58507
rect 10067 58448 10123 58504
rect 10920 58452 10976 58508
rect 11088 58451 11144 58507
rect 15667 58448 15723 58504
rect 16520 58452 16576 58508
rect 16688 58451 16744 58507
rect 21267 58448 21323 58504
rect 22120 58452 22176 58508
rect 22288 58451 22344 58507
rect 26867 58448 26923 58504
rect 27720 58452 27776 58508
rect 27888 58451 27944 58507
rect 32467 58448 32523 58504
rect 33320 58452 33376 58508
rect 33488 58451 33544 58507
rect 38067 58448 38123 58504
rect 38920 58452 38976 58508
rect 39088 58451 39144 58507
rect 43667 58448 43723 58504
rect 1667 57122 1723 57178
rect 7267 57122 7323 57178
rect 12867 57122 12923 57178
rect 18467 57122 18523 57178
rect 24067 57122 24123 57178
rect 29667 57122 29723 57178
rect 35267 57122 35323 57178
rect 40867 57122 40923 57178
rect 448 56896 504 56952
rect 6048 56896 6104 56952
rect 11648 56896 11704 56952
rect 17248 56896 17304 56952
rect 22848 56896 22904 56952
rect 28448 56896 28504 56952
rect 34048 56896 34104 56952
rect 39648 56896 39704 56952
rect 4435 56504 4491 56560
rect 10035 56504 10091 56560
rect 15635 56504 15691 56560
rect 21235 56504 21291 56560
rect 26835 56504 26891 56560
rect 32435 56504 32491 56560
rect 38035 56504 38091 56560
rect 43635 56504 43691 56560
rect 44128 56504 44184 56560
rect -280 56168 -224 56224
rect 1344 56168 1400 56224
rect 5320 56168 5376 56224
rect 6944 56168 7000 56224
rect 10920 56168 10976 56224
rect 12544 56168 12600 56224
rect 16520 56168 16576 56224
rect 18144 56168 18200 56224
rect 22120 56168 22176 56224
rect 23744 56168 23800 56224
rect 27720 56168 27776 56224
rect 29344 56168 29400 56224
rect 33320 56168 33376 56224
rect 34944 56168 35000 56224
rect 38920 56168 38976 56224
rect 40544 56168 40600 56224
rect -112 55776 -56 55832
rect 5488 55776 5544 55832
rect 11088 55776 11144 55832
rect 16688 55776 16744 55832
rect 22288 55776 22344 55832
rect 27888 55776 27944 55832
rect 33488 55776 33544 55832
rect 39088 55776 39144 55832
rect 4467 55440 4523 55496
rect 10067 55440 10123 55496
rect 15667 55440 15723 55496
rect 21267 55440 21323 55496
rect 26867 55440 26923 55496
rect 32467 55440 32523 55496
rect 38067 55440 38123 55496
rect 43667 55440 43723 55496
rect 44128 55440 44184 55496
rect -280 54868 -224 54924
rect -112 54867 -56 54923
rect 4467 54864 4523 54920
rect 5320 54868 5376 54924
rect 5488 54867 5544 54923
rect 10067 54864 10123 54920
rect 10920 54868 10976 54924
rect 11088 54867 11144 54923
rect 15667 54864 15723 54920
rect 16520 54868 16576 54924
rect 16688 54867 16744 54923
rect 21267 54864 21323 54920
rect 22120 54868 22176 54924
rect 22288 54867 22344 54923
rect 26867 54864 26923 54920
rect 27720 54868 27776 54924
rect 27888 54867 27944 54923
rect 32467 54864 32523 54920
rect 33320 54868 33376 54924
rect 33488 54867 33544 54923
rect 38067 54864 38123 54920
rect 38920 54868 38976 54924
rect 39088 54867 39144 54923
rect 43667 54864 43723 54920
rect 1667 53538 1723 53594
rect 7267 53538 7323 53594
rect 12867 53538 12923 53594
rect 18467 53538 18523 53594
rect 24067 53538 24123 53594
rect 29667 53538 29723 53594
rect 35267 53538 35323 53594
rect 40867 53538 40923 53594
rect 448 53312 504 53368
rect 6048 53312 6104 53368
rect 11648 53312 11704 53368
rect 17248 53312 17304 53368
rect 22848 53312 22904 53368
rect 28448 53312 28504 53368
rect 34048 53312 34104 53368
rect 39648 53312 39704 53368
rect 4435 52920 4491 52976
rect 10035 52920 10091 52976
rect 15635 52920 15691 52976
rect 21235 52920 21291 52976
rect 26835 52920 26891 52976
rect 32435 52920 32491 52976
rect 38035 52920 38091 52976
rect 43635 52920 43691 52976
rect 44128 52920 44184 52976
rect -280 52584 -224 52640
rect 1344 52584 1400 52640
rect 5320 52584 5376 52640
rect 6944 52584 7000 52640
rect 10920 52584 10976 52640
rect 12544 52584 12600 52640
rect 16520 52584 16576 52640
rect 18144 52584 18200 52640
rect 22120 52584 22176 52640
rect 23744 52584 23800 52640
rect 27720 52584 27776 52640
rect 29344 52584 29400 52640
rect 33320 52584 33376 52640
rect 34944 52584 35000 52640
rect 38920 52584 38976 52640
rect 40544 52584 40600 52640
rect -112 52192 -56 52248
rect 5488 52192 5544 52248
rect 11088 52192 11144 52248
rect 16688 52192 16744 52248
rect 22288 52192 22344 52248
rect 27888 52192 27944 52248
rect 33488 52192 33544 52248
rect 39088 52192 39144 52248
rect 4467 51856 4523 51912
rect 10067 51856 10123 51912
rect 15667 51856 15723 51912
rect 21267 51856 21323 51912
rect 26867 51856 26923 51912
rect 32467 51856 32523 51912
rect 38067 51856 38123 51912
rect 43667 51856 43723 51912
rect 44128 51856 44184 51912
rect -280 51284 -224 51340
rect -112 51283 -56 51339
rect 4467 51280 4523 51336
rect 5320 51284 5376 51340
rect 5488 51283 5544 51339
rect 10067 51280 10123 51336
rect 10920 51284 10976 51340
rect 11088 51283 11144 51339
rect 15667 51280 15723 51336
rect 16520 51284 16576 51340
rect 16688 51283 16744 51339
rect 21267 51280 21323 51336
rect 22120 51284 22176 51340
rect 22288 51283 22344 51339
rect 26867 51280 26923 51336
rect 27720 51284 27776 51340
rect 27888 51283 27944 51339
rect 32467 51280 32523 51336
rect 33320 51284 33376 51340
rect 33488 51283 33544 51339
rect 38067 51280 38123 51336
rect 38920 51284 38976 51340
rect 39088 51283 39144 51339
rect 43667 51280 43723 51336
rect 1667 49954 1723 50010
rect 7267 49954 7323 50010
rect 12867 49954 12923 50010
rect 18467 49954 18523 50010
rect 24067 49954 24123 50010
rect 29667 49954 29723 50010
rect 35267 49954 35323 50010
rect 40867 49954 40923 50010
rect 448 49728 504 49784
rect 6048 49728 6104 49784
rect 11648 49728 11704 49784
rect 17248 49728 17304 49784
rect 22848 49728 22904 49784
rect 28448 49728 28504 49784
rect 34048 49728 34104 49784
rect 39648 49728 39704 49784
rect 4435 49336 4491 49392
rect 10035 49336 10091 49392
rect 15635 49336 15691 49392
rect 21235 49336 21291 49392
rect 26835 49336 26891 49392
rect 32435 49336 32491 49392
rect 38035 49336 38091 49392
rect 43635 49336 43691 49392
rect 44128 49336 44184 49392
rect -280 49000 -224 49056
rect 1344 49000 1400 49056
rect 5320 49000 5376 49056
rect 6944 49000 7000 49056
rect 10920 49000 10976 49056
rect 12544 49000 12600 49056
rect 16520 49000 16576 49056
rect 18144 49000 18200 49056
rect 22120 49000 22176 49056
rect 23744 49000 23800 49056
rect 27720 49000 27776 49056
rect 29344 49000 29400 49056
rect 33320 49000 33376 49056
rect 34944 49000 35000 49056
rect 38920 49000 38976 49056
rect 40544 49000 40600 49056
rect -112 48608 -56 48664
rect 5488 48608 5544 48664
rect 11088 48608 11144 48664
rect 16688 48608 16744 48664
rect 22288 48608 22344 48664
rect 27888 48608 27944 48664
rect 33488 48608 33544 48664
rect 39088 48608 39144 48664
rect 4467 48272 4523 48328
rect 10067 48272 10123 48328
rect 15667 48272 15723 48328
rect 21267 48272 21323 48328
rect 26867 48272 26923 48328
rect 32467 48272 32523 48328
rect 38067 48272 38123 48328
rect 43667 48272 43723 48328
rect 44128 48272 44184 48328
rect -280 47699 -224 47755
rect -112 47699 -56 47755
rect 4467 47696 4523 47752
rect 5320 47700 5376 47756
rect 5488 47699 5544 47755
rect 10067 47696 10123 47752
rect 10920 47700 10976 47756
rect 11088 47699 11144 47755
rect 15667 47696 15723 47752
rect 16520 47699 16576 47755
rect 16688 47699 16744 47755
rect 21267 47696 21323 47752
rect 22120 47700 22176 47756
rect 22288 47699 22344 47755
rect 26867 47696 26923 47752
rect 27720 47700 27776 47756
rect 27888 47699 27944 47755
rect 32467 47696 32523 47752
rect 33320 47700 33376 47756
rect 33488 47699 33544 47755
rect 38067 47696 38123 47752
rect 38920 47700 38976 47756
rect 39088 47699 39144 47755
rect 43667 47696 43723 47752
rect 1667 46370 1723 46426
rect 7267 46370 7323 46426
rect 12867 46370 12923 46426
rect 18467 46370 18523 46426
rect 24067 46370 24123 46426
rect 29667 46370 29723 46426
rect 35267 46370 35323 46426
rect 40867 46370 40923 46426
rect 448 46144 504 46200
rect 6048 46144 6104 46200
rect 11648 46144 11704 46200
rect 17248 46144 17304 46200
rect 22848 46144 22904 46200
rect 28448 46144 28504 46200
rect 34048 46144 34104 46200
rect 39648 46144 39704 46200
rect 4435 45752 4491 45808
rect 10035 45752 10091 45808
rect 15635 45752 15691 45808
rect 21235 45752 21291 45808
rect 26835 45752 26891 45808
rect 32435 45752 32491 45808
rect 38035 45752 38091 45808
rect 43635 45752 43691 45808
rect 44128 45752 44184 45808
rect -280 45416 -224 45472
rect 1344 45416 1400 45472
rect 5320 45416 5376 45472
rect 6944 45416 7000 45472
rect 10920 45416 10976 45472
rect 12544 45416 12600 45472
rect 16520 45416 16576 45472
rect 18144 45416 18200 45472
rect 22120 45416 22176 45472
rect 23744 45416 23800 45472
rect 27720 45416 27776 45472
rect 29344 45416 29400 45472
rect 33320 45416 33376 45472
rect 34944 45416 35000 45472
rect 38920 45416 38976 45472
rect 40544 45416 40600 45472
rect -112 45024 -56 45080
rect 5488 45024 5544 45080
rect 11088 45024 11144 45080
rect 16688 45024 16744 45080
rect 22288 45024 22344 45080
rect 27888 45024 27944 45080
rect 33488 45024 33544 45080
rect 39088 45024 39144 45080
rect 4467 44688 4523 44744
rect 10067 44688 10123 44744
rect 15667 44688 15723 44744
rect 21267 44688 21323 44744
rect 26867 44688 26923 44744
rect 32467 44688 32523 44744
rect 38067 44688 38123 44744
rect 43667 44688 43723 44744
rect 44128 44688 44184 44744
rect -280 44116 -224 44172
rect -112 44115 -56 44171
rect 4467 44112 4523 44168
rect 5320 44116 5376 44172
rect 5488 44115 5544 44171
rect 10067 44112 10123 44168
rect 10920 44116 10976 44172
rect 11088 44115 11144 44171
rect 15667 44112 15723 44168
rect 16520 44116 16576 44172
rect 16688 44115 16744 44171
rect 21267 44112 21323 44168
rect 22120 44116 22176 44172
rect 22288 44115 22344 44171
rect 26867 44112 26923 44168
rect 27720 44116 27776 44172
rect 27888 44115 27944 44171
rect 32467 44112 32523 44168
rect 33320 44116 33376 44172
rect 33488 44115 33544 44171
rect 38067 44112 38123 44168
rect 38920 44116 38976 44172
rect 39088 44115 39144 44171
rect 43667 44116 43723 44172
rect 2264 42784 2320 42840
rect 7864 42784 7920 42840
rect 13463 42784 13519 42840
rect 19064 42784 19120 42840
rect 24663 42784 24719 42840
rect 30263 42784 30319 42840
rect 35863 42784 35919 42840
rect 41463 42784 41519 42840
rect 448 42560 504 42616
rect 6048 42560 6104 42616
rect 11648 42560 11704 42616
rect 17248 42560 17304 42616
rect 22848 42560 22904 42616
rect 28448 42560 28504 42616
rect 34048 42560 34104 42616
rect 39648 42560 39704 42616
rect 4435 42168 4491 42224
rect 10035 42168 10091 42224
rect 15635 42168 15691 42224
rect 21235 42168 21291 42224
rect 26835 42168 26891 42224
rect 32435 42168 32491 42224
rect 38035 42168 38091 42224
rect 43635 42168 43691 42224
rect 44128 42168 44184 42224
rect 45024 69776 45136 69832
rect 45024 66192 45136 66248
rect 45024 62608 45136 62664
rect 45024 59024 45136 59080
rect 45024 55440 45136 55496
rect 45024 51856 45136 51912
rect 45024 48272 45136 48328
rect 45024 44688 45136 44744
rect 45499 67256 45611 67312
rect 45497 63672 45609 63728
rect 45499 60088 45611 60144
rect 45497 56504 45609 56560
rect 45498 52920 45610 52976
rect 45500 49336 45612 49392
rect 45497 45752 45609 45808
rect 45498 42168 45610 42224
<< metal2 >>
rect -616 67704 -448 70461
rect -122 70168 -46 70179
rect -122 70112 -112 70168
rect -56 70112 -46 70168
rect -122 70103 -46 70112
rect -112 69269 -56 70103
rect 4456 69832 4532 69843
rect 4456 69776 4467 69832
rect 4523 69776 4532 69832
rect 4456 69767 4532 69776
rect -122 69259 -46 69269
rect 4467 69265 4523 69767
rect -122 69203 -112 69259
rect -56 69203 -46 69259
rect -122 69193 -46 69203
rect 4456 69256 4532 69265
rect 4456 69200 4467 69256
rect 4523 69200 4532 69256
rect 4456 69189 4532 69200
rect 1650 67930 1750 67934
rect 1344 67874 1667 67930
rect 1723 67874 1750 67930
rect 439 67704 515 67715
rect -616 67648 448 67704
rect 504 67648 515 67704
rect -616 64120 -448 67648
rect 439 67639 515 67648
rect 1344 66986 1400 67874
rect 1650 67870 1750 67874
rect 4435 67324 4491 68146
rect 4984 67704 5152 70460
rect 5478 70168 5554 70179
rect 5478 70112 5488 70168
rect 5544 70112 5554 70168
rect 5478 70103 5554 70112
rect 5488 69269 5544 70103
rect 10056 69832 10132 69843
rect 10056 69776 10067 69832
rect 10123 69776 10132 69832
rect 10056 69767 10132 69776
rect 5478 69259 5554 69269
rect 10067 69265 10123 69767
rect 5478 69203 5488 69259
rect 5544 69203 5554 69259
rect 5478 69193 5554 69203
rect 10056 69256 10132 69265
rect 10056 69200 10067 69256
rect 10123 69200 10132 69256
rect 10056 69189 10132 69200
rect 7250 67930 7350 67934
rect 6944 67874 7267 67930
rect 7323 67874 7350 67930
rect 6039 67704 6115 67715
rect 4984 67648 6048 67704
rect 6104 67648 6115 67704
rect 4424 67312 4500 67324
rect 4424 67256 4435 67312
rect 4491 67256 4500 67312
rect 4424 67248 4500 67256
rect -290 66976 -214 66986
rect -290 66920 -280 66976
rect -224 66920 -214 66976
rect -290 66910 -214 66920
rect 1335 66976 1411 66986
rect 1335 66920 1344 66976
rect 1400 66920 1411 66976
rect 1335 66910 1411 66920
rect -280 65688 -224 66910
rect -122 66584 -46 66595
rect -122 66528 -112 66584
rect -56 66528 -46 66584
rect -122 66519 -46 66528
rect -290 65676 -214 65688
rect -112 65685 -56 66519
rect 4456 66248 4532 66259
rect 4456 66192 4467 66248
rect 4523 66192 4532 66248
rect 4456 66183 4532 66192
rect -290 65620 -280 65676
rect -224 65620 -214 65676
rect -290 65612 -214 65620
rect -122 65675 -46 65685
rect 4467 65681 4523 66183
rect -122 65619 -112 65675
rect -56 65619 -46 65675
rect -122 65609 -46 65619
rect 4456 65672 4532 65681
rect 4456 65616 4467 65672
rect 4523 65616 4532 65672
rect 4456 65605 4532 65616
rect 1650 64346 1750 64350
rect 1344 64290 1667 64346
rect 1723 64290 1750 64346
rect 439 64120 515 64131
rect -616 64064 448 64120
rect 504 64064 515 64120
rect -616 60536 -448 64064
rect 439 64055 515 64064
rect -290 63392 -214 63403
rect 1344 63402 1400 64290
rect 1650 64286 1750 64290
rect 4435 63740 4491 64562
rect 4984 64120 5152 67648
rect 6039 67639 6115 67648
rect 5310 66976 5386 66987
rect 6944 66986 7000 67874
rect 7250 67870 7350 67874
rect 10035 67324 10091 68146
rect 10584 67704 10752 70516
rect 11078 70168 11154 70179
rect 11078 70112 11088 70168
rect 11144 70112 11154 70168
rect 11078 70103 11154 70112
rect 11088 69269 11144 70103
rect 15656 69832 15732 69843
rect 15656 69776 15667 69832
rect 15723 69776 15732 69832
rect 15656 69767 15732 69776
rect 11078 69259 11154 69269
rect 15667 69265 15723 69767
rect 11078 69203 11088 69259
rect 11144 69203 11154 69259
rect 11078 69193 11154 69203
rect 15656 69256 15732 69265
rect 15656 69200 15667 69256
rect 15723 69200 15732 69256
rect 15656 69189 15732 69200
rect 12850 67930 12950 67934
rect 12544 67874 12867 67930
rect 12923 67874 12950 67930
rect 11639 67704 11715 67715
rect 10584 67648 11648 67704
rect 11704 67648 11715 67704
rect 10024 67312 10100 67324
rect 10024 67256 10035 67312
rect 10091 67256 10100 67312
rect 10024 67248 10100 67256
rect 5310 66920 5320 66976
rect 5376 66920 5386 66976
rect 5310 66911 5386 66920
rect 6935 66976 7011 66986
rect 6935 66920 6944 66976
rect 7000 66920 7011 66976
rect 5320 65688 5376 66911
rect 6935 66910 7011 66920
rect 5478 66584 5554 66595
rect 5478 66528 5488 66584
rect 5544 66528 5554 66584
rect 5478 66519 5554 66528
rect 5310 65676 5386 65688
rect 5488 65685 5544 66519
rect 10056 66248 10132 66259
rect 10056 66192 10067 66248
rect 10123 66192 10132 66248
rect 10056 66183 10132 66192
rect 5310 65620 5320 65676
rect 5376 65620 5386 65676
rect 5310 65612 5386 65620
rect 5478 65675 5554 65685
rect 10067 65681 10123 66183
rect 5478 65619 5488 65675
rect 5544 65619 5554 65675
rect 5478 65609 5554 65619
rect 10056 65672 10132 65681
rect 10056 65616 10067 65672
rect 10123 65616 10132 65672
rect 10056 65605 10132 65616
rect 7250 64346 7350 64350
rect 6944 64290 7267 64346
rect 7323 64290 7350 64346
rect 6039 64120 6115 64131
rect 4984 64064 6048 64120
rect 6104 64064 6115 64120
rect 4424 63728 4500 63740
rect 4424 63672 4435 63728
rect 4491 63672 4500 63728
rect 4424 63664 4500 63672
rect -290 63336 -280 63392
rect -224 63336 -214 63392
rect -290 63327 -214 63336
rect 1335 63392 1411 63402
rect 1335 63336 1344 63392
rect 1400 63336 1411 63392
rect -280 62104 -224 63327
rect 1335 63326 1411 63336
rect -122 63000 -46 63011
rect -122 62944 -112 63000
rect -56 62944 -46 63000
rect -122 62935 -46 62944
rect -290 62092 -214 62104
rect -112 62101 -56 62935
rect 4456 62664 4532 62675
rect 4456 62608 4467 62664
rect 4523 62608 4532 62664
rect 4456 62599 4532 62608
rect -290 62036 -280 62092
rect -224 62036 -214 62092
rect -290 62028 -214 62036
rect -122 62091 -46 62101
rect 4467 62097 4523 62599
rect -122 62035 -112 62091
rect -56 62035 -46 62091
rect -122 62025 -46 62035
rect 4456 62088 4532 62097
rect 4456 62032 4467 62088
rect 4523 62032 4532 62088
rect 4456 62021 4532 62032
rect 1650 60762 1750 60766
rect 1344 60706 1667 60762
rect 1723 60706 1750 60762
rect 439 60536 515 60547
rect -616 60480 448 60536
rect 504 60480 515 60536
rect -616 56952 -448 60480
rect 439 60471 515 60480
rect -290 59808 -214 59820
rect 1344 59818 1400 60706
rect 1650 60702 1750 60706
rect 4435 60156 4491 60978
rect 4984 60536 5152 64064
rect 6039 64055 6115 64064
rect 5310 63392 5386 63404
rect 6944 63402 7000 64290
rect 7250 64286 7350 64290
rect 10035 63740 10091 64562
rect 10584 64120 10752 67648
rect 11639 67639 11715 67648
rect 10910 66976 10986 66987
rect 12544 66986 12600 67874
rect 12850 67870 12950 67874
rect 15635 67324 15691 68146
rect 16184 67704 16352 70461
rect 16678 70168 16754 70179
rect 16678 70112 16688 70168
rect 16744 70112 16754 70168
rect 16678 70103 16754 70112
rect 16688 69269 16744 70103
rect 21256 69832 21332 69843
rect 21256 69776 21267 69832
rect 21323 69776 21332 69832
rect 21256 69767 21332 69776
rect 16678 69259 16754 69269
rect 21267 69265 21323 69767
rect 16678 69203 16688 69259
rect 16744 69203 16754 69259
rect 16678 69193 16754 69203
rect 21256 69256 21332 69265
rect 21256 69200 21267 69256
rect 21323 69200 21332 69256
rect 21256 69189 21332 69200
rect 18450 67930 18550 67934
rect 18144 67874 18467 67930
rect 18523 67874 18550 67930
rect 17239 67704 17315 67715
rect 16184 67648 17248 67704
rect 17304 67648 17315 67704
rect 15624 67312 15700 67324
rect 15624 67256 15635 67312
rect 15691 67256 15700 67312
rect 15624 67248 15700 67256
rect 10910 66920 10920 66976
rect 10976 66920 10986 66976
rect 10910 66911 10986 66920
rect 12535 66976 12611 66986
rect 12535 66920 12544 66976
rect 12600 66920 12611 66976
rect 10920 65688 10976 66911
rect 12535 66910 12611 66920
rect 11078 66584 11154 66595
rect 11078 66528 11088 66584
rect 11144 66528 11154 66584
rect 11078 66519 11154 66528
rect 10910 65676 10986 65688
rect 11088 65685 11144 66519
rect 15656 66248 15732 66259
rect 15656 66192 15667 66248
rect 15723 66192 15732 66248
rect 15656 66183 15732 66192
rect 10910 65620 10920 65676
rect 10976 65620 10986 65676
rect 10910 65612 10986 65620
rect 11078 65675 11154 65685
rect 15667 65681 15723 66183
rect 11078 65619 11088 65675
rect 11144 65619 11154 65675
rect 11078 65609 11154 65619
rect 15656 65672 15732 65681
rect 15656 65616 15667 65672
rect 15723 65616 15732 65672
rect 15656 65605 15732 65616
rect 12850 64346 12950 64350
rect 12544 64290 12867 64346
rect 12923 64290 12950 64346
rect 11639 64120 11715 64131
rect 10584 64064 11648 64120
rect 11704 64064 11715 64120
rect 10024 63728 10100 63740
rect 10024 63672 10035 63728
rect 10091 63672 10100 63728
rect 10024 63664 10100 63672
rect 5310 63336 5320 63392
rect 5376 63336 5386 63392
rect 5310 63328 5386 63336
rect 6935 63392 7011 63402
rect 6935 63336 6944 63392
rect 7000 63336 7011 63392
rect 5320 62104 5376 63328
rect 6935 63326 7011 63336
rect 5478 63000 5554 63011
rect 5478 62944 5488 63000
rect 5544 62944 5554 63000
rect 5478 62935 5554 62944
rect 5310 62092 5386 62104
rect 5488 62101 5544 62935
rect 10056 62664 10132 62675
rect 10056 62608 10067 62664
rect 10123 62608 10132 62664
rect 10056 62599 10132 62608
rect 5310 62036 5320 62092
rect 5376 62036 5386 62092
rect 5310 62028 5386 62036
rect 5478 62091 5554 62101
rect 10067 62097 10123 62599
rect 5478 62035 5488 62091
rect 5544 62035 5554 62091
rect 5478 62025 5554 62035
rect 10056 62088 10132 62097
rect 10056 62032 10067 62088
rect 10123 62032 10132 62088
rect 10056 62021 10132 62032
rect 7250 60762 7350 60766
rect 6944 60706 7267 60762
rect 7323 60706 7350 60762
rect 6039 60536 6115 60547
rect 4984 60480 6048 60536
rect 6104 60480 6115 60536
rect 4424 60144 4500 60156
rect 4424 60088 4435 60144
rect 4491 60088 4500 60144
rect 4424 60080 4500 60088
rect -290 59752 -280 59808
rect -224 59752 -214 59808
rect -290 59744 -214 59752
rect 1335 59808 1411 59818
rect 1335 59752 1344 59808
rect 1400 59752 1411 59808
rect -280 58520 -224 59744
rect 1335 59742 1411 59752
rect -122 59416 -46 59427
rect -122 59360 -112 59416
rect -56 59360 -46 59416
rect -122 59351 -46 59360
rect -290 58508 -214 58520
rect -112 58517 -56 59351
rect 4456 59080 4532 59091
rect 4456 59024 4467 59080
rect 4523 59024 4532 59080
rect 4456 59015 4532 59024
rect -290 58452 -280 58508
rect -224 58452 -214 58508
rect -290 58444 -214 58452
rect -122 58507 -46 58517
rect 4467 58513 4523 59015
rect -122 58451 -112 58507
rect -56 58451 -46 58507
rect -122 58441 -46 58451
rect 4456 58504 4532 58513
rect 4456 58448 4467 58504
rect 4523 58448 4532 58504
rect 4456 58437 4532 58448
rect 1650 57178 1750 57182
rect 1344 57122 1667 57178
rect 1723 57122 1750 57178
rect 439 56952 515 56963
rect -616 56896 448 56952
rect 504 56896 515 56952
rect -616 53368 -448 56896
rect 439 56887 515 56896
rect -289 56224 -213 56235
rect 1344 56234 1400 57122
rect 1650 57118 1750 57122
rect 4435 56572 4491 57394
rect 4984 56952 5152 60480
rect 6039 60471 6115 60480
rect 5310 59808 5386 59819
rect 6944 59818 7000 60706
rect 7250 60702 7350 60706
rect 10035 60156 10091 60978
rect 10584 60536 10752 64064
rect 11639 64055 11715 64064
rect 10910 63392 10986 63403
rect 12544 63402 12600 64290
rect 12850 64286 12950 64290
rect 15635 63740 15691 64562
rect 16184 64120 16352 67648
rect 17239 67639 17315 67648
rect 16511 66976 16587 66987
rect 18144 66986 18200 67874
rect 18450 67870 18550 67874
rect 21235 67324 21291 68146
rect 21784 67704 21952 70459
rect 22278 70168 22354 70179
rect 22278 70112 22288 70168
rect 22344 70112 22354 70168
rect 22278 70103 22354 70112
rect 22288 69269 22344 70103
rect 26856 69832 26932 69843
rect 26856 69776 26867 69832
rect 26923 69776 26932 69832
rect 26856 69767 26932 69776
rect 22278 69259 22354 69269
rect 26867 69265 26923 69767
rect 22278 69203 22288 69259
rect 22344 69203 22354 69259
rect 22278 69193 22354 69203
rect 26856 69256 26932 69265
rect 26856 69200 26867 69256
rect 26923 69200 26932 69256
rect 26856 69189 26932 69200
rect 24050 67930 24150 67934
rect 23744 67874 24067 67930
rect 24123 67874 24150 67930
rect 22839 67704 22915 67715
rect 21784 67648 22848 67704
rect 22904 67648 22915 67704
rect 21224 67312 21300 67324
rect 21224 67256 21235 67312
rect 21291 67256 21300 67312
rect 21224 67248 21300 67256
rect 16511 66920 16520 66976
rect 16576 66920 16587 66976
rect 16511 66911 16587 66920
rect 18135 66976 18211 66986
rect 18135 66920 18144 66976
rect 18200 66920 18211 66976
rect 16520 65688 16576 66911
rect 18135 66910 18211 66920
rect 16678 66584 16754 66595
rect 16678 66528 16688 66584
rect 16744 66528 16754 66584
rect 16678 66519 16754 66528
rect 16510 65676 16586 65688
rect 16688 65685 16744 66519
rect 21256 66248 21332 66259
rect 21256 66192 21267 66248
rect 21323 66192 21332 66248
rect 21256 66183 21332 66192
rect 16510 65620 16520 65676
rect 16576 65620 16586 65676
rect 16510 65612 16586 65620
rect 16678 65675 16754 65685
rect 21267 65681 21323 66183
rect 16678 65619 16688 65675
rect 16744 65619 16754 65675
rect 16678 65609 16754 65619
rect 21256 65672 21332 65681
rect 21256 65616 21267 65672
rect 21323 65616 21332 65672
rect 21256 65605 21332 65616
rect 18450 64346 18550 64350
rect 18144 64290 18467 64346
rect 18523 64290 18550 64346
rect 17239 64120 17315 64131
rect 16184 64064 17248 64120
rect 17304 64064 17315 64120
rect 15624 63728 15700 63740
rect 15624 63672 15635 63728
rect 15691 63672 15700 63728
rect 15624 63664 15700 63672
rect 10910 63336 10920 63392
rect 10976 63336 10986 63392
rect 10910 63327 10986 63336
rect 12535 63392 12611 63402
rect 12535 63336 12544 63392
rect 12600 63336 12611 63392
rect 10920 62104 10976 63327
rect 12535 63326 12611 63336
rect 11078 63000 11154 63011
rect 11078 62944 11088 63000
rect 11144 62944 11154 63000
rect 11078 62935 11154 62944
rect 10910 62092 10986 62104
rect 11088 62101 11144 62935
rect 15656 62664 15732 62675
rect 15656 62608 15667 62664
rect 15723 62608 15732 62664
rect 15656 62599 15732 62608
rect 10910 62036 10920 62092
rect 10976 62036 10986 62092
rect 10910 62028 10986 62036
rect 11078 62091 11154 62101
rect 15667 62097 15723 62599
rect 11078 62035 11088 62091
rect 11144 62035 11154 62091
rect 11078 62025 11154 62035
rect 15656 62088 15732 62097
rect 15656 62032 15667 62088
rect 15723 62032 15732 62088
rect 15656 62021 15732 62032
rect 12850 60762 12950 60766
rect 12544 60706 12867 60762
rect 12923 60706 12950 60762
rect 11639 60536 11715 60547
rect 10584 60480 11648 60536
rect 11704 60480 11715 60536
rect 10024 60144 10100 60156
rect 10024 60088 10035 60144
rect 10091 60088 10100 60144
rect 10024 60080 10100 60088
rect 5310 59752 5320 59808
rect 5376 59752 5386 59808
rect 5310 59743 5386 59752
rect 6935 59808 7011 59818
rect 6935 59752 6944 59808
rect 7000 59752 7011 59808
rect 5320 58520 5376 59743
rect 6935 59742 7011 59752
rect 5478 59416 5554 59427
rect 5478 59360 5488 59416
rect 5544 59360 5554 59416
rect 5478 59351 5554 59360
rect 5310 58508 5386 58520
rect 5488 58517 5544 59351
rect 10056 59080 10132 59091
rect 10056 59024 10067 59080
rect 10123 59024 10132 59080
rect 10056 59015 10132 59024
rect 5310 58452 5320 58508
rect 5376 58452 5386 58508
rect 5310 58444 5386 58452
rect 5478 58507 5554 58517
rect 10067 58513 10123 59015
rect 5478 58451 5488 58507
rect 5544 58451 5554 58507
rect 5478 58441 5554 58451
rect 10056 58504 10132 58513
rect 10056 58448 10067 58504
rect 10123 58448 10132 58504
rect 10056 58437 10132 58448
rect 7250 57178 7350 57182
rect 6944 57122 7267 57178
rect 7323 57122 7350 57178
rect 6039 56952 6115 56963
rect 4984 56896 6048 56952
rect 6104 56896 6115 56952
rect 4424 56560 4500 56572
rect 4424 56504 4435 56560
rect 4491 56504 4500 56560
rect 4424 56496 4500 56504
rect -289 56168 -280 56224
rect -224 56168 -213 56224
rect -289 56159 -213 56168
rect 1335 56224 1411 56234
rect 1335 56168 1344 56224
rect 1400 56168 1411 56224
rect -280 54936 -224 56159
rect 1335 56158 1411 56168
rect -122 55832 -46 55843
rect -122 55776 -112 55832
rect -56 55776 -46 55832
rect -122 55767 -46 55776
rect -290 54924 -214 54936
rect -112 54933 -56 55767
rect 4456 55496 4532 55507
rect 4456 55440 4467 55496
rect 4523 55440 4532 55496
rect 4456 55431 4532 55440
rect -290 54868 -280 54924
rect -224 54868 -214 54924
rect -290 54860 -214 54868
rect -122 54923 -46 54933
rect 4467 54929 4523 55431
rect -122 54867 -112 54923
rect -56 54867 -46 54923
rect -122 54857 -46 54867
rect 4456 54920 4532 54929
rect 4456 54864 4467 54920
rect 4523 54864 4532 54920
rect 4456 54853 4532 54864
rect 1650 53594 1750 53598
rect 1344 53538 1667 53594
rect 1723 53538 1750 53594
rect 439 53368 515 53379
rect -616 53312 448 53368
rect 504 53312 515 53368
rect -616 49784 -448 53312
rect 439 53303 515 53312
rect -290 52640 -214 52651
rect 1344 52650 1400 53538
rect 1650 53534 1750 53538
rect 4435 52988 4491 53810
rect 4984 53368 5152 56896
rect 6039 56887 6115 56896
rect 5310 56224 5386 56236
rect 6944 56234 7000 57122
rect 7250 57118 7350 57122
rect 10035 56572 10091 57394
rect 10584 56952 10752 60480
rect 11639 60471 11715 60480
rect 10910 59808 10986 59819
rect 12544 59818 12600 60706
rect 12850 60702 12950 60706
rect 15635 60156 15691 60978
rect 16184 60536 16352 64064
rect 17239 64055 17315 64064
rect 16511 63392 16587 63404
rect 18144 63402 18200 64290
rect 18450 64286 18550 64290
rect 21235 63740 21291 64562
rect 21784 64120 21952 67648
rect 22839 67639 22915 67648
rect 23744 66986 23800 67874
rect 24050 67870 24150 67874
rect 26835 67324 26891 68146
rect 27384 67704 27552 70478
rect 27878 70168 27954 70179
rect 27878 70112 27888 70168
rect 27944 70112 27954 70168
rect 27878 70103 27954 70112
rect 27888 69269 27944 70103
rect 32456 69832 32532 69843
rect 32456 69776 32467 69832
rect 32523 69776 32532 69832
rect 32456 69767 32532 69776
rect 27878 69259 27954 69269
rect 32467 69265 32523 69767
rect 27878 69203 27888 69259
rect 27944 69203 27954 69259
rect 27878 69193 27954 69203
rect 32456 69256 32532 69265
rect 32456 69200 32467 69256
rect 32523 69200 32532 69256
rect 32456 69189 32532 69200
rect 29650 67930 29750 67934
rect 29344 67874 29667 67930
rect 29723 67874 29750 67930
rect 28439 67704 28515 67715
rect 27384 67648 28448 67704
rect 28504 67648 28515 67704
rect 26824 67312 26900 67324
rect 26824 67256 26835 67312
rect 26891 67256 26900 67312
rect 26824 67248 26900 67256
rect 22110 66976 22186 66986
rect 22110 66920 22120 66976
rect 22176 66920 22186 66976
rect 22110 66910 22186 66920
rect 23735 66976 23811 66986
rect 23735 66920 23744 66976
rect 23800 66920 23811 66976
rect 23735 66910 23811 66920
rect 22120 65688 22176 66910
rect 22278 66584 22354 66595
rect 22278 66528 22288 66584
rect 22344 66528 22354 66584
rect 22278 66519 22354 66528
rect 22110 65676 22186 65688
rect 22288 65685 22344 66519
rect 26856 66248 26932 66259
rect 26856 66192 26867 66248
rect 26923 66192 26932 66248
rect 26856 66183 26932 66192
rect 22110 65620 22120 65676
rect 22176 65620 22186 65676
rect 22110 65612 22186 65620
rect 22278 65675 22354 65685
rect 26867 65681 26923 66183
rect 22278 65619 22288 65675
rect 22344 65619 22354 65675
rect 22278 65609 22354 65619
rect 26856 65672 26932 65681
rect 26856 65616 26867 65672
rect 26923 65616 26932 65672
rect 26856 65605 26932 65616
rect 24050 64346 24150 64350
rect 23744 64290 24067 64346
rect 24123 64290 24150 64346
rect 22839 64120 22915 64131
rect 21784 64064 22848 64120
rect 22904 64064 22915 64120
rect 21224 63728 21300 63740
rect 21224 63672 21235 63728
rect 21291 63672 21300 63728
rect 21224 63664 21300 63672
rect 16511 63336 16520 63392
rect 16576 63336 16587 63392
rect 16511 63328 16587 63336
rect 18135 63392 18211 63402
rect 18135 63336 18144 63392
rect 18200 63336 18211 63392
rect 16520 62104 16576 63328
rect 18135 63326 18211 63336
rect 16678 63000 16754 63011
rect 16678 62944 16688 63000
rect 16744 62944 16754 63000
rect 16678 62935 16754 62944
rect 16510 62092 16586 62104
rect 16688 62101 16744 62935
rect 21256 62664 21332 62675
rect 21256 62608 21267 62664
rect 21323 62608 21332 62664
rect 21256 62599 21332 62608
rect 16510 62036 16520 62092
rect 16576 62036 16586 62092
rect 16510 62028 16586 62036
rect 16678 62091 16754 62101
rect 21267 62097 21323 62599
rect 16678 62035 16688 62091
rect 16744 62035 16754 62091
rect 16678 62025 16754 62035
rect 21256 62088 21332 62097
rect 21256 62032 21267 62088
rect 21323 62032 21332 62088
rect 21256 62021 21332 62032
rect 18450 60762 18550 60766
rect 18144 60706 18467 60762
rect 18523 60706 18550 60762
rect 17239 60536 17315 60547
rect 16184 60480 17248 60536
rect 17304 60480 17315 60536
rect 15624 60144 15700 60156
rect 15624 60088 15635 60144
rect 15691 60088 15700 60144
rect 15624 60080 15700 60088
rect 10910 59752 10920 59808
rect 10976 59752 10986 59808
rect 10910 59743 10986 59752
rect 12535 59808 12611 59818
rect 12535 59752 12544 59808
rect 12600 59752 12611 59808
rect 10920 58520 10976 59743
rect 12535 59742 12611 59752
rect 11078 59416 11154 59427
rect 11078 59360 11088 59416
rect 11144 59360 11154 59416
rect 11078 59351 11154 59360
rect 10910 58508 10986 58520
rect 11088 58517 11144 59351
rect 15656 59080 15732 59091
rect 15656 59024 15667 59080
rect 15723 59024 15732 59080
rect 15656 59015 15732 59024
rect 10910 58452 10920 58508
rect 10976 58452 10986 58508
rect 10910 58444 10986 58452
rect 11078 58507 11154 58517
rect 15667 58513 15723 59015
rect 11078 58451 11088 58507
rect 11144 58451 11154 58507
rect 11078 58441 11154 58451
rect 15656 58504 15732 58513
rect 15656 58448 15667 58504
rect 15723 58448 15732 58504
rect 15656 58437 15732 58448
rect 12850 57178 12950 57182
rect 12544 57122 12867 57178
rect 12923 57122 12950 57178
rect 11639 56952 11715 56963
rect 10584 56896 11648 56952
rect 11704 56896 11715 56952
rect 10024 56560 10100 56572
rect 10024 56504 10035 56560
rect 10091 56504 10100 56560
rect 10024 56496 10100 56504
rect 5310 56168 5320 56224
rect 5376 56168 5386 56224
rect 5310 56160 5386 56168
rect 6935 56224 7011 56234
rect 6935 56168 6944 56224
rect 7000 56168 7011 56224
rect 5320 54936 5376 56160
rect 6935 56158 7011 56168
rect 5478 55832 5554 55843
rect 5478 55776 5488 55832
rect 5544 55776 5554 55832
rect 5478 55767 5554 55776
rect 5309 54924 5385 54936
rect 5488 54933 5544 55767
rect 10056 55496 10132 55507
rect 10056 55440 10067 55496
rect 10123 55440 10132 55496
rect 10056 55431 10132 55440
rect 5309 54868 5320 54924
rect 5376 54868 5385 54924
rect 5309 54860 5385 54868
rect 5478 54923 5554 54933
rect 10067 54929 10123 55431
rect 5478 54867 5488 54923
rect 5544 54867 5554 54923
rect 5478 54857 5554 54867
rect 10056 54920 10132 54929
rect 10056 54864 10067 54920
rect 10123 54864 10132 54920
rect 10056 54853 10132 54864
rect 7250 53594 7350 53598
rect 6944 53538 7267 53594
rect 7323 53538 7350 53594
rect 6039 53368 6115 53379
rect 4984 53312 6048 53368
rect 6104 53312 6115 53368
rect 4424 52976 4500 52988
rect 4424 52920 4435 52976
rect 4491 52920 4500 52976
rect 4424 52912 4500 52920
rect -290 52584 -280 52640
rect -224 52584 -214 52640
rect -290 52575 -214 52584
rect 1335 52640 1411 52650
rect 1335 52584 1344 52640
rect 1400 52584 1411 52640
rect -280 51352 -224 52575
rect 1335 52574 1411 52584
rect -122 52248 -46 52259
rect -122 52192 -112 52248
rect -56 52192 -46 52248
rect -122 52183 -46 52192
rect -291 51340 -215 51352
rect -112 51349 -56 52183
rect 4456 51912 4532 51923
rect 4456 51856 4467 51912
rect 4523 51856 4532 51912
rect 4456 51847 4532 51856
rect -291 51284 -280 51340
rect -224 51284 -215 51340
rect -291 51276 -215 51284
rect -122 51339 -46 51349
rect 4467 51345 4523 51847
rect -122 51283 -112 51339
rect -56 51283 -46 51339
rect -122 51273 -46 51283
rect 4456 51336 4532 51345
rect 4456 51280 4467 51336
rect 4523 51280 4532 51336
rect 4456 51269 4532 51280
rect 1650 50010 1750 50014
rect 1344 49954 1667 50010
rect 1723 49954 1750 50010
rect 439 49784 515 49795
rect -616 49728 448 49784
rect 504 49728 515 49784
rect -616 46200 -448 49728
rect 439 49719 515 49728
rect -290 49056 -214 49067
rect 1344 49066 1400 49954
rect 1650 49950 1750 49954
rect 4435 49404 4491 50226
rect 4984 49784 5152 53312
rect 6039 53303 6115 53312
rect 5310 52640 5386 52651
rect 6944 52650 7000 53538
rect 7250 53534 7350 53538
rect 10035 52988 10091 53810
rect 10584 53368 10752 56896
rect 11639 56887 11715 56896
rect 10910 56224 10986 56235
rect 12544 56234 12600 57122
rect 12850 57118 12950 57122
rect 15635 56572 15691 57394
rect 16184 56952 16352 60480
rect 17239 60471 17315 60480
rect 18144 59818 18200 60706
rect 18450 60702 18550 60706
rect 21235 60156 21291 60978
rect 21784 60536 21952 64064
rect 22839 64055 22915 64064
rect 23744 63402 23800 64290
rect 24050 64286 24150 64290
rect 26835 63740 26891 64562
rect 27384 64120 27552 67648
rect 28439 67639 28515 67648
rect 27710 66976 27786 66987
rect 29344 66986 29400 67874
rect 29650 67870 29750 67874
rect 32435 67324 32491 68146
rect 32984 67704 33152 70467
rect 33478 70168 33554 70179
rect 33478 70112 33488 70168
rect 33544 70112 33554 70168
rect 33478 70103 33554 70112
rect 33488 69269 33544 70103
rect 38056 69832 38132 69843
rect 38056 69776 38067 69832
rect 38123 69776 38132 69832
rect 38056 69767 38132 69776
rect 44072 69832 45192 69888
rect 44072 69776 44128 69832
rect 44184 69776 45024 69832
rect 45136 69776 45192 69832
rect 33478 69259 33554 69269
rect 38067 69265 38123 69767
rect 44072 69720 45192 69776
rect 33478 69203 33488 69259
rect 33544 69203 33554 69259
rect 33478 69193 33554 69203
rect 38056 69256 38132 69265
rect 38056 69200 38067 69256
rect 38123 69200 38132 69256
rect 38056 69189 38132 69200
rect 35250 67930 35350 67934
rect 34944 67874 35267 67930
rect 35323 67874 35350 67930
rect 34039 67704 34115 67715
rect 32984 67648 34048 67704
rect 34104 67648 34115 67704
rect 32424 67312 32500 67324
rect 32424 67256 32435 67312
rect 32491 67256 32500 67312
rect 32424 67248 32500 67256
rect 27710 66920 27720 66976
rect 27776 66920 27786 66976
rect 27710 66911 27786 66920
rect 29335 66976 29411 66986
rect 29335 66920 29344 66976
rect 29400 66920 29411 66976
rect 27720 65688 27776 66911
rect 29335 66910 29411 66920
rect 27878 66584 27954 66595
rect 27878 66528 27888 66584
rect 27944 66528 27954 66584
rect 27878 66519 27954 66528
rect 27710 65676 27786 65688
rect 27888 65685 27944 66519
rect 32456 66248 32532 66259
rect 32456 66192 32467 66248
rect 32523 66192 32532 66248
rect 32456 66183 32532 66192
rect 27710 65620 27720 65676
rect 27776 65620 27786 65676
rect 27710 65612 27786 65620
rect 27878 65675 27954 65685
rect 32467 65681 32523 66183
rect 27878 65619 27888 65675
rect 27944 65619 27954 65675
rect 27878 65609 27954 65619
rect 32456 65672 32532 65681
rect 32456 65616 32467 65672
rect 32523 65616 32532 65672
rect 32456 65605 32532 65616
rect 29650 64346 29750 64350
rect 29344 64290 29667 64346
rect 29723 64290 29750 64346
rect 28439 64120 28515 64131
rect 27384 64064 28448 64120
rect 28504 64064 28515 64120
rect 26824 63728 26900 63740
rect 26824 63672 26835 63728
rect 26891 63672 26900 63728
rect 26824 63664 26900 63672
rect 22110 63392 22186 63402
rect 22110 63336 22120 63392
rect 22176 63336 22186 63392
rect 22110 63326 22186 63336
rect 23735 63392 23811 63402
rect 23735 63336 23744 63392
rect 23800 63336 23811 63392
rect 23735 63326 23811 63336
rect 22120 62104 22176 63326
rect 22278 63000 22354 63011
rect 22278 62944 22288 63000
rect 22344 62944 22354 63000
rect 22278 62935 22354 62944
rect 22110 62092 22186 62104
rect 22288 62101 22344 62935
rect 26856 62664 26932 62675
rect 26856 62608 26867 62664
rect 26923 62608 26932 62664
rect 26856 62599 26932 62608
rect 22110 62036 22120 62092
rect 22176 62036 22186 62092
rect 22110 62028 22186 62036
rect 22278 62091 22354 62101
rect 26867 62097 26923 62599
rect 22278 62035 22288 62091
rect 22344 62035 22354 62091
rect 22278 62025 22354 62035
rect 26856 62088 26932 62097
rect 26856 62032 26867 62088
rect 26923 62032 26932 62088
rect 26856 62021 26932 62032
rect 24050 60762 24150 60766
rect 23744 60706 24067 60762
rect 24123 60706 24150 60762
rect 22839 60536 22915 60547
rect 21784 60480 22848 60536
rect 22904 60480 22915 60536
rect 21224 60144 21300 60156
rect 21224 60088 21235 60144
rect 21291 60088 21300 60144
rect 21224 60080 21300 60088
rect 16509 59808 16585 59818
rect 16509 59752 16520 59808
rect 16576 59752 16585 59808
rect 16509 59742 16585 59752
rect 18135 59808 18211 59818
rect 18135 59752 18144 59808
rect 18200 59752 18211 59808
rect 18135 59742 18211 59752
rect 16520 58520 16576 59742
rect 16678 59416 16754 59427
rect 16678 59360 16688 59416
rect 16744 59360 16754 59416
rect 16678 59351 16754 59360
rect 16510 58508 16586 58520
rect 16688 58517 16744 59351
rect 21256 59080 21332 59091
rect 21256 59024 21267 59080
rect 21323 59024 21332 59080
rect 21256 59015 21332 59024
rect 16510 58452 16520 58508
rect 16576 58452 16586 58508
rect 16510 58444 16586 58452
rect 16678 58507 16754 58517
rect 21267 58513 21323 59015
rect 16678 58451 16688 58507
rect 16744 58451 16754 58507
rect 16678 58441 16754 58451
rect 21256 58504 21332 58513
rect 21256 58448 21267 58504
rect 21323 58448 21332 58504
rect 21256 58437 21332 58448
rect 18450 57178 18550 57182
rect 18144 57122 18467 57178
rect 18523 57122 18550 57178
rect 17239 56952 17315 56963
rect 16184 56896 17248 56952
rect 17304 56896 17315 56952
rect 15624 56560 15700 56572
rect 15624 56504 15635 56560
rect 15691 56504 15700 56560
rect 15624 56496 15700 56504
rect 10910 56168 10920 56224
rect 10976 56168 10986 56224
rect 10910 56159 10986 56168
rect 12535 56224 12611 56234
rect 12535 56168 12544 56224
rect 12600 56168 12611 56224
rect 10920 54936 10976 56159
rect 12535 56158 12611 56168
rect 11078 55832 11154 55843
rect 11078 55776 11088 55832
rect 11144 55776 11154 55832
rect 11078 55767 11154 55776
rect 10910 54924 10986 54936
rect 11088 54933 11144 55767
rect 15656 55496 15732 55507
rect 15656 55440 15667 55496
rect 15723 55440 15732 55496
rect 15656 55431 15732 55440
rect 10910 54868 10920 54924
rect 10976 54868 10986 54924
rect 10910 54860 10986 54868
rect 11078 54923 11154 54933
rect 15667 54929 15723 55431
rect 11078 54867 11088 54923
rect 11144 54867 11154 54923
rect 11078 54857 11154 54867
rect 15656 54920 15732 54929
rect 15656 54864 15667 54920
rect 15723 54864 15732 54920
rect 15656 54853 15732 54864
rect 12850 53594 12950 53598
rect 12544 53538 12867 53594
rect 12923 53538 12950 53594
rect 11639 53368 11715 53379
rect 10584 53312 11648 53368
rect 11704 53312 11715 53368
rect 10024 52976 10100 52988
rect 10024 52920 10035 52976
rect 10091 52920 10100 52976
rect 10024 52912 10100 52920
rect 5310 52584 5320 52640
rect 5376 52584 5386 52640
rect 5310 52575 5386 52584
rect 6935 52640 7011 52650
rect 6935 52584 6944 52640
rect 7000 52584 7011 52640
rect 5320 51352 5376 52575
rect 6935 52574 7011 52584
rect 5478 52248 5554 52259
rect 5478 52192 5488 52248
rect 5544 52192 5554 52248
rect 5478 52183 5554 52192
rect 5310 51340 5386 51352
rect 5488 51349 5544 52183
rect 10056 51912 10132 51923
rect 10056 51856 10067 51912
rect 10123 51856 10132 51912
rect 10056 51847 10132 51856
rect 5310 51284 5320 51340
rect 5376 51284 5386 51340
rect 5310 51276 5386 51284
rect 5478 51339 5554 51349
rect 10067 51345 10123 51847
rect 5478 51283 5488 51339
rect 5544 51283 5554 51339
rect 5478 51273 5554 51283
rect 10056 51336 10132 51345
rect 10056 51280 10067 51336
rect 10123 51280 10132 51336
rect 10056 51269 10132 51280
rect 7250 50010 7350 50014
rect 6944 49954 7267 50010
rect 7323 49954 7350 50010
rect 6039 49784 6115 49795
rect 4984 49728 6048 49784
rect 6104 49728 6115 49784
rect 4424 49392 4500 49404
rect 4424 49336 4435 49392
rect 4491 49336 4500 49392
rect 4424 49328 4500 49336
rect -290 49000 -280 49056
rect -224 49000 -214 49056
rect -290 48991 -214 49000
rect 1335 49056 1411 49066
rect 1335 49000 1344 49056
rect 1400 49000 1411 49056
rect -280 47766 -224 48991
rect 1335 48990 1411 49000
rect -122 48664 -46 48675
rect -122 48608 -112 48664
rect -56 48608 -46 48664
rect -122 48599 -46 48608
rect -291 47755 -215 47766
rect -112 47765 -56 48599
rect 4456 48328 4532 48339
rect 4456 48272 4467 48328
rect 4523 48272 4532 48328
rect 4456 48263 4532 48272
rect -291 47699 -280 47755
rect -224 47699 -215 47755
rect -291 47690 -215 47699
rect -122 47755 -46 47765
rect 4467 47761 4523 48263
rect -122 47699 -112 47755
rect -56 47699 -46 47755
rect -122 47689 -46 47699
rect 4456 47752 4532 47761
rect 4456 47696 4467 47752
rect 4523 47696 4532 47752
rect 4456 47685 4532 47696
rect 1650 46426 1750 46430
rect 1344 46370 1667 46426
rect 1723 46370 1750 46426
rect 439 46200 515 46211
rect -616 46144 448 46200
rect 504 46144 515 46200
rect -616 42616 -448 46144
rect 439 46135 515 46144
rect -291 45472 -215 45483
rect 1344 45482 1400 46370
rect 1650 46366 1750 46370
rect 4435 45820 4491 46642
rect 4984 46200 5152 49728
rect 6039 49719 6115 49728
rect 5310 49056 5386 49067
rect 6944 49066 7000 49954
rect 7250 49950 7350 49954
rect 10035 49404 10091 50226
rect 10584 49784 10752 53312
rect 11639 53303 11715 53312
rect 10910 52640 10986 52651
rect 12544 52650 12600 53538
rect 12850 53534 12950 53538
rect 15635 52988 15691 53810
rect 16184 53368 16352 56896
rect 17239 56887 17315 56896
rect 16510 56224 16586 56237
rect 18144 56234 18200 57122
rect 18450 57118 18550 57122
rect 21235 56572 21291 57394
rect 21784 56952 21952 60480
rect 22839 60471 22915 60480
rect 22109 59808 22185 59819
rect 23744 59818 23800 60706
rect 24050 60702 24150 60706
rect 26835 60156 26891 60978
rect 27384 60536 27552 64064
rect 28439 64055 28515 64064
rect 27710 63392 27786 63403
rect 29344 63402 29400 64290
rect 29650 64286 29750 64290
rect 32435 63740 32491 64562
rect 32984 64120 33152 67648
rect 34039 67639 34115 67648
rect 33310 66976 33386 66987
rect 34944 66986 35000 67874
rect 35250 67870 35350 67874
rect 38035 67324 38091 68146
rect 38024 67312 38100 67324
rect 38024 67256 38035 67312
rect 38091 67256 38100 67312
rect 38024 67248 38100 67256
rect 33310 66920 33320 66976
rect 33376 66920 33386 66976
rect 33310 66911 33386 66920
rect 34935 66976 35011 66986
rect 34935 66920 34944 66976
rect 35000 66920 35011 66976
rect 33320 65688 33376 66911
rect 34935 66910 35011 66920
rect 33478 66584 33554 66595
rect 33478 66528 33488 66584
rect 33544 66528 33554 66584
rect 33478 66519 33554 66528
rect 33310 65676 33386 65688
rect 33488 65685 33544 66519
rect 38056 66248 38132 66259
rect 38056 66192 38067 66248
rect 38123 66192 38132 66248
rect 38056 66183 38132 66192
rect 33310 65620 33320 65676
rect 33376 65620 33386 65676
rect 33310 65612 33386 65620
rect 33478 65675 33554 65685
rect 38067 65681 38123 66183
rect 33478 65619 33488 65675
rect 33544 65619 33554 65675
rect 33478 65609 33554 65619
rect 38056 65672 38132 65681
rect 38056 65616 38067 65672
rect 38123 65616 38132 65672
rect 38056 65605 38132 65616
rect 35250 64346 35350 64350
rect 34944 64290 35267 64346
rect 35323 64290 35350 64346
rect 34039 64120 34115 64131
rect 32984 64064 34048 64120
rect 34104 64064 34115 64120
rect 32424 63728 32500 63740
rect 32424 63672 32435 63728
rect 32491 63672 32500 63728
rect 32424 63664 32500 63672
rect 27710 63336 27720 63392
rect 27776 63336 27786 63392
rect 27710 63327 27786 63336
rect 29335 63392 29411 63402
rect 29335 63336 29344 63392
rect 29400 63336 29411 63392
rect 27720 62104 27776 63327
rect 29335 63326 29411 63336
rect 27878 63000 27954 63011
rect 27878 62944 27888 63000
rect 27944 62944 27954 63000
rect 27878 62935 27954 62944
rect 27710 62092 27786 62104
rect 27888 62101 27944 62935
rect 32456 62664 32532 62675
rect 32456 62608 32467 62664
rect 32523 62608 32532 62664
rect 32456 62599 32532 62608
rect 27710 62036 27720 62092
rect 27776 62036 27786 62092
rect 27710 62028 27786 62036
rect 27878 62091 27954 62101
rect 32467 62097 32523 62599
rect 27878 62035 27888 62091
rect 27944 62035 27954 62091
rect 27878 62025 27954 62035
rect 32456 62088 32532 62097
rect 32456 62032 32467 62088
rect 32523 62032 32532 62088
rect 32456 62021 32532 62032
rect 29650 60762 29750 60766
rect 29344 60706 29667 60762
rect 29723 60706 29750 60762
rect 28439 60536 28515 60547
rect 27384 60480 28448 60536
rect 28504 60480 28515 60536
rect 26824 60144 26900 60156
rect 26824 60088 26835 60144
rect 26891 60088 26900 60144
rect 26824 60080 26900 60088
rect 22109 59752 22120 59808
rect 22176 59752 22185 59808
rect 22109 59743 22185 59752
rect 23735 59808 23811 59818
rect 23735 59752 23744 59808
rect 23800 59752 23811 59808
rect 22120 58520 22176 59743
rect 23735 59742 23811 59752
rect 22278 59416 22354 59427
rect 22278 59360 22288 59416
rect 22344 59360 22354 59416
rect 22278 59351 22354 59360
rect 22110 58508 22186 58520
rect 22288 58517 22344 59351
rect 26856 59080 26932 59091
rect 26856 59024 26867 59080
rect 26923 59024 26932 59080
rect 26856 59015 26932 59024
rect 22110 58452 22120 58508
rect 22176 58452 22186 58508
rect 22110 58444 22186 58452
rect 22278 58507 22354 58517
rect 26867 58513 26923 59015
rect 22278 58451 22288 58507
rect 22344 58451 22354 58507
rect 22278 58441 22354 58451
rect 26856 58504 26932 58513
rect 26856 58448 26867 58504
rect 26923 58448 26932 58504
rect 26856 58437 26932 58448
rect 24050 57178 24150 57182
rect 23744 57122 24067 57178
rect 24123 57122 24150 57178
rect 22839 56952 22915 56963
rect 21784 56896 22848 56952
rect 22904 56896 22915 56952
rect 21224 56560 21300 56572
rect 21224 56504 21235 56560
rect 21291 56504 21300 56560
rect 21224 56496 21300 56504
rect 16510 56168 16520 56224
rect 16576 56168 16586 56224
rect 16510 56161 16586 56168
rect 18135 56224 18211 56234
rect 18135 56168 18144 56224
rect 18200 56168 18211 56224
rect 16520 54936 16576 56161
rect 18135 56158 18211 56168
rect 16678 55832 16754 55843
rect 16678 55776 16688 55832
rect 16744 55776 16754 55832
rect 16678 55767 16754 55776
rect 16509 54924 16585 54936
rect 16688 54933 16744 55767
rect 21256 55496 21332 55507
rect 21256 55440 21267 55496
rect 21323 55440 21332 55496
rect 21256 55431 21332 55440
rect 16509 54868 16520 54924
rect 16576 54868 16585 54924
rect 16509 54860 16585 54868
rect 16678 54923 16754 54933
rect 21267 54929 21323 55431
rect 16678 54867 16688 54923
rect 16744 54867 16754 54923
rect 16678 54857 16754 54867
rect 21256 54920 21332 54929
rect 21256 54864 21267 54920
rect 21323 54864 21332 54920
rect 21256 54853 21332 54864
rect 18450 53594 18550 53598
rect 18144 53538 18467 53594
rect 18523 53538 18550 53594
rect 17239 53368 17315 53379
rect 16184 53312 17248 53368
rect 17304 53312 17315 53368
rect 15624 52976 15700 52988
rect 15624 52920 15635 52976
rect 15691 52920 15700 52976
rect 15624 52912 15700 52920
rect 10910 52584 10920 52640
rect 10976 52584 10986 52640
rect 10910 52575 10986 52584
rect 12535 52640 12611 52650
rect 12535 52584 12544 52640
rect 12600 52584 12611 52640
rect 10920 51352 10976 52575
rect 12535 52574 12611 52584
rect 11078 52248 11154 52259
rect 11078 52192 11088 52248
rect 11144 52192 11154 52248
rect 11078 52183 11154 52192
rect 10910 51340 10986 51352
rect 11088 51349 11144 52183
rect 15656 51912 15732 51923
rect 15656 51856 15667 51912
rect 15723 51856 15732 51912
rect 15656 51847 15732 51856
rect 10910 51284 10920 51340
rect 10976 51284 10986 51340
rect 10910 51276 10986 51284
rect 11078 51339 11154 51349
rect 15667 51345 15723 51847
rect 11078 51283 11088 51339
rect 11144 51283 11154 51339
rect 11078 51273 11154 51283
rect 15656 51336 15732 51345
rect 15656 51280 15667 51336
rect 15723 51280 15732 51336
rect 15656 51269 15732 51280
rect 12850 50010 12950 50014
rect 12544 49954 12867 50010
rect 12923 49954 12950 50010
rect 11639 49784 11715 49795
rect 10584 49728 11648 49784
rect 11704 49728 11715 49784
rect 10024 49392 10100 49404
rect 10024 49336 10035 49392
rect 10091 49336 10100 49392
rect 10024 49328 10100 49336
rect 5310 49000 5320 49056
rect 5376 49000 5386 49056
rect 5310 48991 5386 49000
rect 6935 49056 7011 49066
rect 6935 49000 6944 49056
rect 7000 49000 7011 49056
rect 5320 47768 5376 48991
rect 6935 48990 7011 49000
rect 5478 48664 5554 48675
rect 5478 48608 5488 48664
rect 5544 48608 5554 48664
rect 5478 48599 5554 48608
rect 5309 47756 5385 47768
rect 5488 47765 5544 48599
rect 10056 48328 10132 48339
rect 10056 48272 10067 48328
rect 10123 48272 10132 48328
rect 10056 48263 10132 48272
rect 5309 47700 5320 47756
rect 5376 47700 5385 47756
rect 5309 47692 5385 47700
rect 5478 47755 5554 47765
rect 10067 47761 10123 48263
rect 5478 47699 5488 47755
rect 5544 47699 5554 47755
rect 5478 47689 5554 47699
rect 10056 47752 10132 47761
rect 10056 47696 10067 47752
rect 10123 47696 10132 47752
rect 10056 47685 10132 47696
rect 7250 46426 7350 46430
rect 6944 46370 7267 46426
rect 7323 46370 7350 46426
rect 6039 46200 6115 46211
rect 4984 46144 6048 46200
rect 6104 46144 6115 46200
rect 4424 45808 4500 45820
rect 4424 45752 4435 45808
rect 4491 45752 4500 45808
rect 4424 45744 4500 45752
rect -291 45416 -280 45472
rect -224 45416 -215 45472
rect -291 45407 -215 45416
rect 1335 45472 1411 45482
rect 1335 45416 1344 45472
rect 1400 45416 1411 45472
rect -280 44184 -224 45407
rect 1335 45406 1411 45416
rect -122 45080 -46 45091
rect -122 45024 -112 45080
rect -56 45024 -46 45080
rect -122 45015 -46 45024
rect -290 44172 -214 44184
rect -112 44181 -56 45015
rect 4456 44744 4532 44755
rect 4456 44688 4467 44744
rect 4523 44688 4532 44744
rect 4456 44679 4532 44688
rect -290 44116 -280 44172
rect -224 44116 -214 44172
rect -290 44108 -214 44116
rect -122 44171 -46 44181
rect 4467 44177 4523 44679
rect -122 44115 -112 44171
rect -56 44115 -46 44171
rect -122 44105 -46 44115
rect 4456 44168 4532 44177
rect 4456 44112 4467 44168
rect 4523 44112 4532 44168
rect 4456 44101 4532 44112
rect 2255 42840 2331 42851
rect 2255 42784 2264 42840
rect 2320 42784 2688 42840
rect 2744 42784 2800 42840
rect 2255 42775 2331 42784
rect 439 42616 515 42627
rect -616 42560 448 42616
rect 504 42560 515 42616
rect -616 41776 -448 42560
rect 439 42551 515 42560
rect 4435 42236 4491 43058
rect 4984 42616 5152 46144
rect 6039 46135 6115 46144
rect 5310 45472 5386 45483
rect 6944 45482 7000 46370
rect 7250 46366 7350 46370
rect 10035 45820 10091 46642
rect 10584 46200 10752 49728
rect 11639 49719 11715 49728
rect 12544 49066 12600 49954
rect 12850 49950 12950 49954
rect 15635 49404 15691 50226
rect 16184 49784 16352 53312
rect 17239 53303 17315 53312
rect 18144 52650 18200 53538
rect 18450 53534 18550 53538
rect 21235 52988 21291 53810
rect 21784 53368 21952 56896
rect 22839 56887 22915 56896
rect 22110 56224 22186 56235
rect 23744 56234 23800 57122
rect 24050 57118 24150 57122
rect 26835 56572 26891 57394
rect 27384 56952 27552 60480
rect 28439 60471 28515 60480
rect 29344 59818 29400 60706
rect 29650 60702 29750 60706
rect 32435 60156 32491 60978
rect 32984 60536 33152 64064
rect 34039 64055 34115 64064
rect 33310 63392 33386 63403
rect 34944 63402 35000 64290
rect 35250 64286 35350 64290
rect 38035 63740 38091 64562
rect 38584 64120 38752 69419
rect 44072 67312 45696 67368
rect 44072 67256 44128 67312
rect 44184 67256 45499 67312
rect 45611 67256 45696 67312
rect 44072 67200 45696 67256
rect 38910 66976 38986 66987
rect 38910 66920 38920 66976
rect 38976 66920 38986 66976
rect 38910 66911 38986 66920
rect 38920 65688 38976 66911
rect 39078 66584 39154 66595
rect 39078 66528 39088 66584
rect 39144 66528 39154 66584
rect 39078 66519 39154 66528
rect 38910 65676 38986 65688
rect 39088 65685 39144 66519
rect 43656 66248 43732 66259
rect 43656 66192 43667 66248
rect 43723 66192 43732 66248
rect 43656 66183 43732 66192
rect 44072 66248 45192 66304
rect 44072 66192 44128 66248
rect 44184 66192 45024 66248
rect 45136 66192 45192 66248
rect 38910 65620 38920 65676
rect 38976 65620 38986 65676
rect 38910 65612 38986 65620
rect 39078 65675 39154 65685
rect 43667 65681 43723 66183
rect 44072 66136 45192 66192
rect 39078 65619 39088 65675
rect 39144 65619 39154 65675
rect 39078 65609 39154 65619
rect 43656 65672 43732 65681
rect 43656 65616 43667 65672
rect 43723 65616 43732 65672
rect 43656 65605 43732 65616
rect 40850 64346 40950 64350
rect 40544 64290 40867 64346
rect 40923 64290 40950 64346
rect 39639 64120 39715 64131
rect 38584 64064 39648 64120
rect 39704 64064 39715 64120
rect 38024 63728 38100 63740
rect 38024 63672 38035 63728
rect 38091 63672 38100 63728
rect 38024 63664 38100 63672
rect 33310 63336 33320 63392
rect 33376 63336 33386 63392
rect 33310 63327 33386 63336
rect 34935 63392 35011 63402
rect 34935 63336 34944 63392
rect 35000 63336 35011 63392
rect 33320 62104 33376 63327
rect 34935 63326 35011 63336
rect 33478 63000 33554 63011
rect 33478 62944 33488 63000
rect 33544 62944 33554 63000
rect 33478 62935 33554 62944
rect 33310 62092 33386 62104
rect 33488 62101 33544 62935
rect 38056 62664 38132 62675
rect 38056 62608 38067 62664
rect 38123 62608 38132 62664
rect 38056 62599 38132 62608
rect 33310 62036 33320 62092
rect 33376 62036 33386 62092
rect 33310 62028 33386 62036
rect 33478 62091 33554 62101
rect 38067 62097 38123 62599
rect 33478 62035 33488 62091
rect 33544 62035 33554 62091
rect 33478 62025 33554 62035
rect 38056 62088 38132 62097
rect 38056 62032 38067 62088
rect 38123 62032 38132 62088
rect 38056 62021 38132 62032
rect 35250 60762 35350 60766
rect 34944 60706 35267 60762
rect 35323 60706 35350 60762
rect 34039 60536 34115 60547
rect 32984 60480 34048 60536
rect 34104 60480 34115 60536
rect 32424 60144 32500 60156
rect 32424 60088 32435 60144
rect 32491 60088 32500 60144
rect 32424 60080 32500 60088
rect 27710 59808 27786 59818
rect 27710 59752 27720 59808
rect 27776 59752 27786 59808
rect 27710 59742 27786 59752
rect 29335 59808 29411 59818
rect 29335 59752 29344 59808
rect 29400 59752 29411 59808
rect 29335 59742 29411 59752
rect 27720 58520 27776 59742
rect 27878 59416 27954 59427
rect 27878 59360 27888 59416
rect 27944 59360 27954 59416
rect 27878 59351 27954 59360
rect 27710 58508 27786 58520
rect 27888 58517 27944 59351
rect 32456 59080 32532 59091
rect 32456 59024 32467 59080
rect 32523 59024 32532 59080
rect 32456 59015 32532 59024
rect 27710 58452 27720 58508
rect 27776 58452 27786 58508
rect 27710 58444 27786 58452
rect 27878 58507 27954 58517
rect 32467 58513 32523 59015
rect 27878 58451 27888 58507
rect 27944 58451 27954 58507
rect 27878 58441 27954 58451
rect 32456 58504 32532 58513
rect 32456 58448 32467 58504
rect 32523 58448 32532 58504
rect 32456 58437 32532 58448
rect 29650 57178 29750 57182
rect 29344 57122 29667 57178
rect 29723 57122 29750 57178
rect 28439 56952 28515 56963
rect 27384 56896 28448 56952
rect 28504 56896 28515 56952
rect 26824 56560 26900 56572
rect 26824 56504 26835 56560
rect 26891 56504 26900 56560
rect 26824 56496 26900 56504
rect 22110 56168 22120 56224
rect 22176 56168 22186 56224
rect 22110 56159 22186 56168
rect 23735 56224 23811 56234
rect 23735 56168 23744 56224
rect 23800 56168 23811 56224
rect 22120 54936 22176 56159
rect 23735 56158 23811 56168
rect 22278 55832 22354 55843
rect 22278 55776 22288 55832
rect 22344 55776 22354 55832
rect 22278 55767 22354 55776
rect 22110 54924 22186 54936
rect 22288 54933 22344 55767
rect 26856 55496 26932 55507
rect 26856 55440 26867 55496
rect 26923 55440 26932 55496
rect 26856 55431 26932 55440
rect 22110 54868 22120 54924
rect 22176 54868 22186 54924
rect 22110 54860 22186 54868
rect 22278 54923 22354 54933
rect 26867 54929 26923 55431
rect 22278 54867 22288 54923
rect 22344 54867 22354 54923
rect 22278 54857 22354 54867
rect 26856 54920 26932 54929
rect 26856 54864 26867 54920
rect 26923 54864 26932 54920
rect 26856 54853 26932 54864
rect 24050 53594 24150 53598
rect 23744 53538 24067 53594
rect 24123 53538 24150 53594
rect 22839 53368 22915 53379
rect 21784 53312 22848 53368
rect 22904 53312 22915 53368
rect 21224 52976 21300 52988
rect 21224 52920 21235 52976
rect 21291 52920 21300 52976
rect 21224 52912 21300 52920
rect 16509 52640 16585 52650
rect 16509 52584 16520 52640
rect 16576 52584 16585 52640
rect 16509 52574 16585 52584
rect 18135 52640 18211 52650
rect 18135 52584 18144 52640
rect 18200 52584 18211 52640
rect 18135 52574 18211 52584
rect 16520 51352 16576 52574
rect 16678 52248 16754 52259
rect 16678 52192 16688 52248
rect 16744 52192 16754 52248
rect 16678 52183 16754 52192
rect 16510 51340 16586 51352
rect 16688 51349 16744 52183
rect 21256 51912 21332 51923
rect 21256 51856 21267 51912
rect 21323 51856 21332 51912
rect 21256 51847 21332 51856
rect 16510 51284 16520 51340
rect 16576 51284 16586 51340
rect 16510 51276 16586 51284
rect 16678 51339 16754 51349
rect 21267 51345 21323 51847
rect 16678 51283 16688 51339
rect 16744 51283 16754 51339
rect 16678 51273 16754 51283
rect 21256 51336 21332 51345
rect 21256 51280 21267 51336
rect 21323 51280 21332 51336
rect 21256 51269 21332 51280
rect 18450 50010 18550 50014
rect 18144 49954 18467 50010
rect 18523 49954 18550 50010
rect 17239 49784 17315 49795
rect 16184 49728 17248 49784
rect 17304 49728 17315 49784
rect 15624 49392 15700 49404
rect 15624 49336 15635 49392
rect 15691 49336 15700 49392
rect 15624 49328 15700 49336
rect 10910 49056 10986 49066
rect 10910 49000 10920 49056
rect 10976 49000 10986 49056
rect 10910 48990 10986 49000
rect 12535 49056 12611 49066
rect 12535 49000 12544 49056
rect 12600 49000 12611 49056
rect 12535 48990 12611 49000
rect 10920 47768 10976 48990
rect 11078 48664 11154 48675
rect 11078 48608 11088 48664
rect 11144 48608 11154 48664
rect 11078 48599 11154 48608
rect 10910 47756 10986 47768
rect 11088 47765 11144 48599
rect 15656 48328 15732 48339
rect 15656 48272 15667 48328
rect 15723 48272 15732 48328
rect 15656 48263 15732 48272
rect 10910 47700 10920 47756
rect 10976 47700 10986 47756
rect 10910 47692 10986 47700
rect 11078 47755 11154 47765
rect 15667 47761 15723 48263
rect 11078 47699 11088 47755
rect 11144 47699 11154 47755
rect 11078 47689 11154 47699
rect 15656 47752 15732 47761
rect 15656 47696 15667 47752
rect 15723 47696 15732 47752
rect 15656 47685 15732 47696
rect 12850 46426 12950 46430
rect 12544 46370 12867 46426
rect 12923 46370 12950 46426
rect 11639 46200 11715 46211
rect 10584 46144 11648 46200
rect 11704 46144 11715 46200
rect 10024 45808 10100 45820
rect 10024 45752 10035 45808
rect 10091 45752 10100 45808
rect 10024 45744 10100 45752
rect 5310 45416 5320 45472
rect 5376 45416 5386 45472
rect 5310 45407 5386 45416
rect 6935 45472 7011 45482
rect 6935 45416 6944 45472
rect 7000 45416 7011 45472
rect 5320 44184 5376 45407
rect 6935 45406 7011 45416
rect 5478 45080 5554 45091
rect 5478 45024 5488 45080
rect 5544 45024 5554 45080
rect 5478 45015 5554 45024
rect 5310 44172 5386 44184
rect 5488 44181 5544 45015
rect 10056 44744 10132 44755
rect 10056 44688 10067 44744
rect 10123 44688 10132 44744
rect 10056 44679 10132 44688
rect 5310 44116 5320 44172
rect 5376 44116 5386 44172
rect 5310 44108 5386 44116
rect 5478 44171 5554 44181
rect 10067 44177 10123 44679
rect 5478 44115 5488 44171
rect 5544 44115 5554 44171
rect 5478 44105 5554 44115
rect 10056 44168 10132 44177
rect 10056 44112 10067 44168
rect 10123 44112 10132 44168
rect 10056 44101 10132 44112
rect 7853 42840 7929 42850
rect 7853 42784 7864 42840
rect 7920 42784 8288 42840
rect 8344 42784 8400 42840
rect 7853 42774 7929 42784
rect 6039 42616 6115 42627
rect 4984 42560 6048 42616
rect 6104 42560 6115 42616
rect 4424 42224 4500 42236
rect 4424 42168 4435 42224
rect 4491 42168 4500 42224
rect 4424 42160 4500 42168
rect 4984 41995 5152 42560
rect 6039 42551 6115 42560
rect 10035 42236 10091 43058
rect 10584 42616 10752 46144
rect 11639 46135 11715 46144
rect 10910 45472 10986 45485
rect 12544 45482 12600 46370
rect 12850 46366 12950 46370
rect 15635 45820 15691 46642
rect 16184 46200 16352 49728
rect 17239 49719 17315 49728
rect 16509 49056 16585 49067
rect 18144 49066 18200 49954
rect 18450 49950 18550 49954
rect 21235 49404 21291 50226
rect 21784 49784 21952 53312
rect 22839 53303 22915 53312
rect 23744 52650 23800 53538
rect 24050 53534 24150 53538
rect 26835 52988 26891 53810
rect 27384 53368 27552 56896
rect 28439 56887 28515 56896
rect 27710 56224 27786 56235
rect 29344 56234 29400 57122
rect 29650 57118 29750 57122
rect 32435 56572 32491 57394
rect 32984 56952 33152 60480
rect 34039 60471 34115 60480
rect 33310 59808 33386 59820
rect 34944 59818 35000 60706
rect 35250 60702 35350 60706
rect 38035 60156 38091 60978
rect 38584 60536 38752 64064
rect 39639 64055 39715 64064
rect 40544 63402 40600 64290
rect 40850 64286 40950 64290
rect 43635 63740 43691 64562
rect 43624 63728 43700 63740
rect 43624 63672 43635 63728
rect 43691 63672 43700 63728
rect 43624 63664 43700 63672
rect 44072 63728 45696 63784
rect 44072 63672 44128 63728
rect 44184 63672 45497 63728
rect 45609 63672 45696 63728
rect 44072 63616 45696 63672
rect 38910 63392 38986 63402
rect 38910 63336 38920 63392
rect 38976 63336 38986 63392
rect 38910 63326 38986 63336
rect 40535 63392 40611 63402
rect 40535 63336 40544 63392
rect 40600 63336 40611 63392
rect 40535 63326 40611 63336
rect 38920 62104 38976 63326
rect 39078 63000 39154 63011
rect 39078 62944 39088 63000
rect 39144 62944 39154 63000
rect 39078 62935 39154 62944
rect 38910 62092 38986 62104
rect 39088 62101 39144 62935
rect 43656 62664 43732 62675
rect 43656 62608 43667 62664
rect 43723 62608 43732 62664
rect 43656 62599 43732 62608
rect 44072 62664 45192 62720
rect 44072 62608 44128 62664
rect 44184 62608 45024 62664
rect 45136 62608 45192 62664
rect 38910 62036 38920 62092
rect 38976 62036 38986 62092
rect 38910 62028 38986 62036
rect 39078 62091 39154 62101
rect 43667 62097 43723 62599
rect 44072 62552 45192 62608
rect 39078 62035 39088 62091
rect 39144 62035 39154 62091
rect 39078 62025 39154 62035
rect 43656 62088 43732 62097
rect 43656 62032 43667 62088
rect 43723 62032 43732 62088
rect 43656 62021 43732 62032
rect 40850 60762 40950 60766
rect 40544 60706 40867 60762
rect 40923 60706 40950 60762
rect 39639 60536 39715 60547
rect 38584 60480 39648 60536
rect 39704 60480 39715 60536
rect 38024 60144 38100 60156
rect 38024 60088 38035 60144
rect 38091 60088 38100 60144
rect 38024 60080 38100 60088
rect 33310 59752 33320 59808
rect 33376 59752 33386 59808
rect 33310 59744 33386 59752
rect 34935 59808 35011 59818
rect 34935 59752 34944 59808
rect 35000 59752 35011 59808
rect 33320 58520 33376 59744
rect 34935 59742 35011 59752
rect 33478 59416 33554 59427
rect 33478 59360 33488 59416
rect 33544 59360 33554 59416
rect 33478 59351 33554 59360
rect 33310 58508 33386 58520
rect 33488 58517 33544 59351
rect 38056 59080 38132 59091
rect 38056 59024 38067 59080
rect 38123 59024 38132 59080
rect 38056 59015 38132 59024
rect 33310 58452 33320 58508
rect 33376 58452 33386 58508
rect 33310 58444 33386 58452
rect 33478 58507 33554 58517
rect 38067 58513 38123 59015
rect 33478 58451 33488 58507
rect 33544 58451 33554 58507
rect 33478 58441 33554 58451
rect 38056 58504 38132 58513
rect 38056 58448 38067 58504
rect 38123 58448 38132 58504
rect 38056 58437 38132 58448
rect 35250 57178 35350 57182
rect 34944 57122 35267 57178
rect 35323 57122 35350 57178
rect 34039 56952 34115 56963
rect 32984 56896 34048 56952
rect 34104 56896 34115 56952
rect 32424 56560 32500 56572
rect 32424 56504 32435 56560
rect 32491 56504 32500 56560
rect 32424 56496 32500 56504
rect 27710 56168 27720 56224
rect 27776 56168 27786 56224
rect 27710 56159 27786 56168
rect 29335 56224 29411 56234
rect 29335 56168 29344 56224
rect 29400 56168 29411 56224
rect 27720 54936 27776 56159
rect 29335 56158 29411 56168
rect 27878 55832 27954 55843
rect 27878 55776 27888 55832
rect 27944 55776 27954 55832
rect 27878 55767 27954 55776
rect 27710 54924 27786 54936
rect 27888 54933 27944 55767
rect 32456 55496 32532 55507
rect 32456 55440 32467 55496
rect 32523 55440 32532 55496
rect 32456 55431 32532 55440
rect 27710 54868 27720 54924
rect 27776 54868 27786 54924
rect 27710 54860 27786 54868
rect 27878 54923 27954 54933
rect 32467 54929 32523 55431
rect 27878 54867 27888 54923
rect 27944 54867 27954 54923
rect 27878 54857 27954 54867
rect 32456 54920 32532 54929
rect 32456 54864 32467 54920
rect 32523 54864 32532 54920
rect 32456 54853 32532 54864
rect 29650 53594 29750 53598
rect 29344 53538 29667 53594
rect 29723 53538 29750 53594
rect 28439 53368 28515 53379
rect 27384 53312 28448 53368
rect 28504 53312 28515 53368
rect 26824 52976 26900 52988
rect 26824 52920 26835 52976
rect 26891 52920 26900 52976
rect 26824 52912 26900 52920
rect 22109 52640 22185 52650
rect 22109 52584 22120 52640
rect 22176 52584 22185 52640
rect 22109 52574 22185 52584
rect 23735 52640 23811 52650
rect 23735 52584 23744 52640
rect 23800 52584 23811 52640
rect 23735 52574 23811 52584
rect 22120 51352 22176 52574
rect 22278 52248 22354 52259
rect 22278 52192 22288 52248
rect 22344 52192 22354 52248
rect 22278 52183 22354 52192
rect 22109 51340 22185 51352
rect 22288 51349 22344 52183
rect 26856 51912 26932 51923
rect 26856 51856 26867 51912
rect 26923 51856 26932 51912
rect 26856 51847 26932 51856
rect 22109 51284 22120 51340
rect 22176 51284 22185 51340
rect 22109 51276 22185 51284
rect 22278 51339 22354 51349
rect 26867 51345 26923 51847
rect 22278 51283 22288 51339
rect 22344 51283 22354 51339
rect 22278 51273 22354 51283
rect 26856 51336 26932 51345
rect 26856 51280 26867 51336
rect 26923 51280 26932 51336
rect 26856 51269 26932 51280
rect 24050 50010 24150 50014
rect 23744 49954 24067 50010
rect 24123 49954 24150 50010
rect 22839 49784 22915 49795
rect 21784 49728 22848 49784
rect 22904 49728 22915 49784
rect 21224 49392 21300 49404
rect 21224 49336 21235 49392
rect 21291 49336 21300 49392
rect 21224 49328 21300 49336
rect 16509 49000 16520 49056
rect 16576 49000 16585 49056
rect 16509 48991 16585 49000
rect 18135 49056 18211 49066
rect 18135 49000 18144 49056
rect 18200 49000 18211 49056
rect 16520 47766 16576 48991
rect 18135 48990 18211 49000
rect 16678 48664 16754 48675
rect 16678 48608 16688 48664
rect 16744 48608 16754 48664
rect 16678 48599 16754 48608
rect 16508 47755 16584 47766
rect 16688 47765 16744 48599
rect 21256 48328 21332 48339
rect 21256 48272 21267 48328
rect 21323 48272 21332 48328
rect 21256 48263 21332 48272
rect 16508 47699 16520 47755
rect 16576 47699 16584 47755
rect 16508 47690 16584 47699
rect 16678 47755 16754 47765
rect 21267 47761 21323 48263
rect 16678 47699 16688 47755
rect 16744 47699 16754 47755
rect 16678 47689 16754 47699
rect 21256 47752 21332 47761
rect 21256 47696 21267 47752
rect 21323 47696 21332 47752
rect 21256 47685 21332 47696
rect 18450 46426 18550 46430
rect 18144 46370 18467 46426
rect 18523 46370 18550 46426
rect 17239 46200 17315 46211
rect 16184 46144 17248 46200
rect 17304 46144 17315 46200
rect 15624 45808 15700 45820
rect 15624 45752 15635 45808
rect 15691 45752 15700 45808
rect 15624 45744 15700 45752
rect 10910 45416 10920 45472
rect 10976 45416 10986 45472
rect 10910 45409 10986 45416
rect 12535 45472 12611 45482
rect 12535 45416 12544 45472
rect 12600 45416 12611 45472
rect 10920 44184 10976 45409
rect 12535 45406 12611 45416
rect 11078 45080 11154 45091
rect 11078 45024 11088 45080
rect 11144 45024 11154 45080
rect 11078 45015 11154 45024
rect 10910 44172 10986 44184
rect 11088 44181 11144 45015
rect 15656 44744 15732 44755
rect 15656 44688 15667 44744
rect 15723 44688 15732 44744
rect 15656 44679 15732 44688
rect 10910 44116 10920 44172
rect 10976 44116 10986 44172
rect 10910 44108 10986 44116
rect 11078 44171 11154 44181
rect 15667 44177 15723 44679
rect 11078 44115 11088 44171
rect 11144 44115 11154 44171
rect 11078 44105 11154 44115
rect 15656 44168 15732 44177
rect 15656 44112 15667 44168
rect 15723 44112 15732 44168
rect 15656 44101 15732 44112
rect 13453 42840 13529 42851
rect 13453 42784 13463 42840
rect 13519 42784 13888 42840
rect 13944 42784 14000 42840
rect 13453 42775 13529 42784
rect 11639 42616 11715 42627
rect 10584 42560 11648 42616
rect 11704 42560 11715 42616
rect 10024 42224 10100 42236
rect 10024 42168 10035 42224
rect 10091 42168 10100 42224
rect 10024 42160 10100 42168
rect 10584 41995 10752 42560
rect 11639 42551 11715 42560
rect 15635 42236 15691 43058
rect 16184 42616 16352 46144
rect 17239 46135 17315 46144
rect 16510 45472 16586 45483
rect 18144 45482 18200 46370
rect 18450 46366 18550 46370
rect 21235 45820 21291 46642
rect 21784 46200 21952 49728
rect 22839 49719 22915 49728
rect 22111 49056 22187 49067
rect 23744 49066 23800 49954
rect 24050 49950 24150 49954
rect 26835 49404 26891 50226
rect 27384 49784 27552 53312
rect 28439 53303 28515 53312
rect 27709 52640 27785 52651
rect 29344 52650 29400 53538
rect 29650 53534 29750 53538
rect 32435 52988 32491 53810
rect 32984 53368 33152 56896
rect 34039 56887 34115 56896
rect 34944 56234 35000 57122
rect 35250 57118 35350 57122
rect 38035 56572 38091 57394
rect 38584 56952 38752 60480
rect 39639 60471 39715 60480
rect 40544 59818 40600 60706
rect 40850 60702 40950 60706
rect 43635 60156 43691 60978
rect 43624 60144 43700 60156
rect 43624 60088 43635 60144
rect 43691 60088 43700 60144
rect 43624 60080 43700 60088
rect 44072 60144 45696 60200
rect 44072 60088 44128 60144
rect 44184 60088 45499 60144
rect 45611 60088 45696 60144
rect 44072 60032 45696 60088
rect 38909 59808 38985 59818
rect 38909 59752 38920 59808
rect 38976 59752 38985 59808
rect 38909 59742 38985 59752
rect 40535 59808 40611 59818
rect 40535 59752 40544 59808
rect 40600 59752 40611 59808
rect 40535 59742 40611 59752
rect 38920 58520 38976 59742
rect 39078 59416 39154 59427
rect 39078 59360 39088 59416
rect 39144 59360 39154 59416
rect 39078 59351 39154 59360
rect 38910 58508 38986 58520
rect 39088 58517 39144 59351
rect 43656 59080 43732 59091
rect 43656 59024 43667 59080
rect 43723 59024 43732 59080
rect 43656 59015 43732 59024
rect 44072 59080 45192 59136
rect 44072 59024 44128 59080
rect 44184 59024 45024 59080
rect 45136 59024 45192 59080
rect 38910 58452 38920 58508
rect 38976 58452 38986 58508
rect 38910 58444 38986 58452
rect 39078 58507 39154 58517
rect 43667 58513 43723 59015
rect 44072 58968 45192 59024
rect 39078 58451 39088 58507
rect 39144 58451 39154 58507
rect 39078 58441 39154 58451
rect 43656 58504 43732 58513
rect 43656 58448 43667 58504
rect 43723 58448 43732 58504
rect 43656 58437 43732 58448
rect 40850 57178 40950 57182
rect 40544 57122 40867 57178
rect 40923 57122 40950 57178
rect 39639 56952 39715 56963
rect 38584 56896 39648 56952
rect 39704 56896 39715 56952
rect 38024 56560 38100 56572
rect 38024 56504 38035 56560
rect 38091 56504 38100 56560
rect 38024 56496 38100 56504
rect 33310 56224 33386 56234
rect 33310 56168 33320 56224
rect 33376 56168 33386 56224
rect 33310 56158 33386 56168
rect 34935 56224 35011 56234
rect 34935 56168 34944 56224
rect 35000 56168 35011 56224
rect 34935 56158 35011 56168
rect 33320 54936 33376 56158
rect 33478 55832 33554 55843
rect 33478 55776 33488 55832
rect 33544 55776 33554 55832
rect 33478 55767 33554 55776
rect 33310 54924 33386 54936
rect 33488 54933 33544 55767
rect 38056 55496 38132 55507
rect 38056 55440 38067 55496
rect 38123 55440 38132 55496
rect 38056 55431 38132 55440
rect 33310 54868 33320 54924
rect 33376 54868 33386 54924
rect 33310 54860 33386 54868
rect 33478 54923 33554 54933
rect 38067 54929 38123 55431
rect 33478 54867 33488 54923
rect 33544 54867 33554 54923
rect 33478 54857 33554 54867
rect 38056 54920 38132 54929
rect 38056 54864 38067 54920
rect 38123 54864 38132 54920
rect 38056 54853 38132 54864
rect 35250 53594 35350 53598
rect 34944 53538 35267 53594
rect 35323 53538 35350 53594
rect 34039 53368 34115 53379
rect 32984 53312 34048 53368
rect 34104 53312 34115 53368
rect 32424 52976 32500 52988
rect 32424 52920 32435 52976
rect 32491 52920 32500 52976
rect 32424 52912 32500 52920
rect 27709 52584 27720 52640
rect 27776 52584 27785 52640
rect 27709 52575 27785 52584
rect 29335 52640 29411 52650
rect 29335 52584 29344 52640
rect 29400 52584 29411 52640
rect 27720 51352 27776 52575
rect 29335 52574 29411 52584
rect 27878 52248 27954 52259
rect 27878 52192 27888 52248
rect 27944 52192 27954 52248
rect 27878 52183 27954 52192
rect 27710 51340 27786 51352
rect 27888 51349 27944 52183
rect 32456 51912 32532 51923
rect 32456 51856 32467 51912
rect 32523 51856 32532 51912
rect 32456 51847 32532 51856
rect 27710 51284 27720 51340
rect 27776 51284 27786 51340
rect 27710 51276 27786 51284
rect 27878 51339 27954 51349
rect 32467 51345 32523 51847
rect 27878 51283 27888 51339
rect 27944 51283 27954 51339
rect 27878 51273 27954 51283
rect 32456 51336 32532 51345
rect 32456 51280 32467 51336
rect 32523 51280 32532 51336
rect 32456 51269 32532 51280
rect 29650 50010 29750 50014
rect 29344 49954 29667 50010
rect 29723 49954 29750 50010
rect 28439 49784 28515 49795
rect 27384 49728 28448 49784
rect 28504 49728 28515 49784
rect 26824 49392 26900 49404
rect 26824 49336 26835 49392
rect 26891 49336 26900 49392
rect 26824 49328 26900 49336
rect 22111 49000 22120 49056
rect 22176 49000 22187 49056
rect 22111 48991 22187 49000
rect 23735 49056 23811 49066
rect 23735 49000 23744 49056
rect 23800 49000 23811 49056
rect 22120 47768 22176 48991
rect 23735 48990 23811 49000
rect 22278 48664 22354 48675
rect 22278 48608 22288 48664
rect 22344 48608 22354 48664
rect 22278 48599 22354 48608
rect 22110 47756 22186 47768
rect 22288 47765 22344 48599
rect 26856 48328 26932 48339
rect 26856 48272 26867 48328
rect 26923 48272 26932 48328
rect 26856 48263 26932 48272
rect 22110 47700 22120 47756
rect 22176 47700 22186 47756
rect 22110 47692 22186 47700
rect 22278 47755 22354 47765
rect 26867 47761 26923 48263
rect 22278 47699 22288 47755
rect 22344 47699 22354 47755
rect 22278 47689 22354 47699
rect 26856 47752 26932 47761
rect 26856 47696 26867 47752
rect 26923 47696 26932 47752
rect 26856 47685 26932 47696
rect 24050 46426 24150 46430
rect 23744 46370 24067 46426
rect 24123 46370 24150 46426
rect 22839 46200 22915 46211
rect 21784 46144 22848 46200
rect 22904 46144 22915 46200
rect 21224 45808 21300 45820
rect 21224 45752 21235 45808
rect 21291 45752 21300 45808
rect 21224 45744 21300 45752
rect 16510 45416 16520 45472
rect 16576 45416 16586 45472
rect 16510 45407 16586 45416
rect 18135 45472 18211 45482
rect 18135 45416 18144 45472
rect 18200 45416 18211 45472
rect 16520 44184 16576 45407
rect 18135 45406 18211 45416
rect 16678 45080 16754 45091
rect 16678 45024 16688 45080
rect 16744 45024 16754 45080
rect 16678 45015 16754 45024
rect 16509 44172 16585 44184
rect 16688 44181 16744 45015
rect 21256 44744 21332 44755
rect 21256 44688 21267 44744
rect 21323 44688 21332 44744
rect 21256 44679 21332 44688
rect 16509 44116 16520 44172
rect 16576 44116 16585 44172
rect 16509 44108 16585 44116
rect 16678 44171 16754 44181
rect 21267 44177 21323 44679
rect 16678 44115 16688 44171
rect 16744 44115 16754 44171
rect 16678 44105 16754 44115
rect 21256 44168 21332 44177
rect 21256 44112 21267 44168
rect 21323 44112 21332 44168
rect 21256 44101 21332 44112
rect 19052 42840 19128 42852
rect 19052 42784 19064 42840
rect 19120 42784 19488 42840
rect 19544 42784 19600 42840
rect 19052 42776 19128 42784
rect 17239 42616 17315 42627
rect 16184 42560 17248 42616
rect 17304 42560 17315 42616
rect 15624 42224 15700 42236
rect 15624 42168 15635 42224
rect 15691 42168 15700 42224
rect 15624 42160 15700 42168
rect 16184 41995 16352 42560
rect 17239 42551 17315 42560
rect 21235 42236 21291 43058
rect 21784 42616 21952 46144
rect 22839 46135 22915 46144
rect 22110 45472 22186 45483
rect 23744 45482 23800 46370
rect 24050 46366 24150 46370
rect 26835 45820 26891 46642
rect 27384 46200 27552 49728
rect 28439 49719 28515 49728
rect 27710 49056 27786 49067
rect 29344 49066 29400 49954
rect 29650 49950 29750 49954
rect 32435 49404 32491 50226
rect 32984 49784 33152 53312
rect 34039 53303 34115 53312
rect 34944 52650 35000 53538
rect 35250 53534 35350 53538
rect 38035 52988 38091 53810
rect 38584 53368 38752 56896
rect 39639 56887 39715 56896
rect 38909 56224 38985 56236
rect 40544 56234 40600 57122
rect 40850 57118 40950 57122
rect 43635 56572 43691 57394
rect 43624 56560 43700 56572
rect 43624 56504 43635 56560
rect 43691 56504 43700 56560
rect 43624 56496 43700 56504
rect 44072 56560 45696 56616
rect 44072 56504 44128 56560
rect 44184 56504 45497 56560
rect 45609 56504 45696 56560
rect 44072 56448 45696 56504
rect 38909 56168 38920 56224
rect 38976 56168 38985 56224
rect 38909 56160 38985 56168
rect 40535 56224 40611 56234
rect 40535 56168 40544 56224
rect 40600 56168 40611 56224
rect 38920 54936 38976 56160
rect 40535 56158 40611 56168
rect 39078 55832 39154 55843
rect 39078 55776 39088 55832
rect 39144 55776 39154 55832
rect 39078 55767 39154 55776
rect 38909 54924 38985 54936
rect 39088 54933 39144 55767
rect 43656 55496 43732 55507
rect 43656 55440 43667 55496
rect 43723 55440 43732 55496
rect 43656 55431 43732 55440
rect 44072 55496 45192 55552
rect 44072 55440 44128 55496
rect 44184 55440 45024 55496
rect 45136 55440 45192 55496
rect 38909 54868 38920 54924
rect 38976 54868 38985 54924
rect 38909 54860 38985 54868
rect 39078 54923 39154 54933
rect 43667 54929 43723 55431
rect 44072 55384 45192 55440
rect 39078 54867 39088 54923
rect 39144 54867 39154 54923
rect 39078 54857 39154 54867
rect 43656 54920 43732 54929
rect 43656 54864 43667 54920
rect 43723 54864 43732 54920
rect 43656 54853 43732 54864
rect 40850 53594 40950 53598
rect 40544 53538 40867 53594
rect 40923 53538 40950 53594
rect 39639 53368 39715 53379
rect 38584 53312 39648 53368
rect 39704 53312 39715 53368
rect 38024 52976 38100 52988
rect 38024 52920 38035 52976
rect 38091 52920 38100 52976
rect 38024 52912 38100 52920
rect 33309 52640 33385 52649
rect 33309 52584 33320 52640
rect 33376 52584 33385 52640
rect 33309 52573 33385 52584
rect 34935 52640 35011 52650
rect 34935 52584 34944 52640
rect 35000 52584 35011 52640
rect 34935 52574 35011 52584
rect 33320 51352 33376 52573
rect 33478 52248 33554 52259
rect 33478 52192 33488 52248
rect 33544 52192 33554 52248
rect 33478 52183 33554 52192
rect 33310 51340 33386 51352
rect 33488 51349 33544 52183
rect 38056 51912 38132 51923
rect 38056 51856 38067 51912
rect 38123 51856 38132 51912
rect 38056 51847 38132 51856
rect 33310 51284 33320 51340
rect 33376 51284 33386 51340
rect 33310 51276 33386 51284
rect 33478 51339 33554 51349
rect 38067 51345 38123 51847
rect 33478 51283 33488 51339
rect 33544 51283 33554 51339
rect 33478 51273 33554 51283
rect 38056 51336 38132 51345
rect 38056 51280 38067 51336
rect 38123 51280 38132 51336
rect 38056 51269 38132 51280
rect 35250 50010 35350 50014
rect 34944 49954 35267 50010
rect 35323 49954 35350 50010
rect 34039 49784 34115 49795
rect 32984 49728 34048 49784
rect 34104 49728 34115 49784
rect 32424 49392 32500 49404
rect 32424 49336 32435 49392
rect 32491 49336 32500 49392
rect 32424 49328 32500 49336
rect 27710 49000 27720 49056
rect 27776 49000 27786 49056
rect 27710 48991 27786 49000
rect 29335 49056 29411 49066
rect 29335 49000 29344 49056
rect 29400 49000 29411 49056
rect 27720 47768 27776 48991
rect 29335 48990 29411 49000
rect 27878 48664 27954 48675
rect 27878 48608 27888 48664
rect 27944 48608 27954 48664
rect 27878 48599 27954 48608
rect 27710 47756 27786 47768
rect 27888 47765 27944 48599
rect 32456 48328 32532 48339
rect 32456 48272 32467 48328
rect 32523 48272 32532 48328
rect 32456 48263 32532 48272
rect 27710 47700 27720 47756
rect 27776 47700 27786 47756
rect 27710 47692 27786 47700
rect 27878 47755 27954 47765
rect 32467 47761 32523 48263
rect 27878 47699 27888 47755
rect 27944 47699 27954 47755
rect 27878 47689 27954 47699
rect 32456 47752 32532 47761
rect 32456 47696 32467 47752
rect 32523 47696 32532 47752
rect 32456 47685 32532 47696
rect 29650 46426 29750 46430
rect 29344 46370 29667 46426
rect 29723 46370 29750 46426
rect 28439 46200 28515 46211
rect 27384 46144 28448 46200
rect 28504 46144 28515 46200
rect 26824 45808 26900 45820
rect 26824 45752 26835 45808
rect 26891 45752 26900 45808
rect 26824 45744 26900 45752
rect 22110 45416 22120 45472
rect 22176 45416 22186 45472
rect 22110 45407 22186 45416
rect 23735 45472 23811 45482
rect 23735 45416 23744 45472
rect 23800 45416 23811 45472
rect 22120 44184 22176 45407
rect 23735 45406 23811 45416
rect 22278 45080 22354 45091
rect 22278 45024 22288 45080
rect 22344 45024 22354 45080
rect 22278 45015 22354 45024
rect 22110 44172 22186 44184
rect 22288 44181 22344 45015
rect 26856 44744 26932 44755
rect 26856 44688 26867 44744
rect 26923 44688 26932 44744
rect 26856 44679 26932 44688
rect 22110 44116 22120 44172
rect 22176 44116 22186 44172
rect 22110 44108 22186 44116
rect 22278 44171 22354 44181
rect 26867 44177 26923 44679
rect 22278 44115 22288 44171
rect 22344 44115 22354 44171
rect 22278 44105 22354 44115
rect 26856 44168 26932 44177
rect 26856 44112 26867 44168
rect 26923 44112 26932 44168
rect 26856 44101 26932 44112
rect 24654 42840 24730 42851
rect 24654 42784 24663 42840
rect 24719 42784 25088 42840
rect 25144 42784 25200 42840
rect 24654 42775 24730 42784
rect 22839 42616 22915 42627
rect 21784 42560 22848 42616
rect 22904 42560 22915 42616
rect 21224 42224 21300 42236
rect 21224 42168 21235 42224
rect 21291 42168 21300 42224
rect 21224 42160 21300 42168
rect 21784 41995 21952 42560
rect 22839 42551 22915 42560
rect 26835 42236 26891 43058
rect 27384 42616 27552 46144
rect 28439 46135 28515 46144
rect 27710 45472 27786 45483
rect 29344 45482 29400 46370
rect 29650 46366 29750 46370
rect 32435 45820 32491 46642
rect 32984 46200 33152 49728
rect 34039 49719 34115 49728
rect 34944 49066 35000 49954
rect 35250 49950 35350 49954
rect 38035 49404 38091 50226
rect 38584 49784 38752 53312
rect 39639 53303 39715 53312
rect 40544 52650 40600 53538
rect 40850 53534 40950 53538
rect 43635 52988 43691 53810
rect 43624 52976 43700 52988
rect 43624 52920 43635 52976
rect 43691 52920 43700 52976
rect 43624 52912 43700 52920
rect 44072 52976 45696 53032
rect 44072 52920 44128 52976
rect 44184 52920 45498 52976
rect 45610 52920 45696 52976
rect 44072 52864 45696 52920
rect 38911 52640 38987 52650
rect 38911 52584 38920 52640
rect 38976 52584 38987 52640
rect 38911 52574 38987 52584
rect 40535 52640 40611 52650
rect 40535 52584 40544 52640
rect 40600 52584 40611 52640
rect 40535 52574 40611 52584
rect 38920 51352 38976 52574
rect 39078 52248 39154 52259
rect 39078 52192 39088 52248
rect 39144 52192 39154 52248
rect 39078 52183 39154 52192
rect 38909 51340 38985 51352
rect 39088 51349 39144 52183
rect 43656 51912 43732 51923
rect 43656 51856 43667 51912
rect 43723 51856 43732 51912
rect 43656 51847 43732 51856
rect 44072 51912 45192 51968
rect 44072 51856 44128 51912
rect 44184 51856 45024 51912
rect 45136 51856 45192 51912
rect 38909 51284 38920 51340
rect 38976 51284 38985 51340
rect 38909 51276 38985 51284
rect 39078 51339 39154 51349
rect 43667 51345 43723 51847
rect 44072 51800 45192 51856
rect 39078 51283 39088 51339
rect 39144 51283 39154 51339
rect 39078 51273 39154 51283
rect 43656 51336 43732 51345
rect 43656 51280 43667 51336
rect 43723 51280 43732 51336
rect 43656 51269 43732 51280
rect 40850 50010 40950 50014
rect 40544 49954 40867 50010
rect 40923 49954 40950 50010
rect 39639 49784 39715 49795
rect 38584 49728 39648 49784
rect 39704 49728 39715 49784
rect 38024 49392 38100 49404
rect 38024 49336 38035 49392
rect 38091 49336 38100 49392
rect 38024 49328 38100 49336
rect 33309 49056 33385 49066
rect 33309 49000 33320 49056
rect 33376 49000 33385 49056
rect 33309 48990 33385 49000
rect 34935 49056 35011 49066
rect 34935 49000 34944 49056
rect 35000 49000 35011 49056
rect 34935 48990 35011 49000
rect 33320 47768 33376 48990
rect 33478 48664 33554 48675
rect 33478 48608 33488 48664
rect 33544 48608 33554 48664
rect 33478 48599 33554 48608
rect 33310 47756 33386 47768
rect 33488 47765 33544 48599
rect 38056 48328 38132 48339
rect 38056 48272 38067 48328
rect 38123 48272 38132 48328
rect 38056 48263 38132 48272
rect 33310 47700 33320 47756
rect 33376 47700 33386 47756
rect 33310 47692 33386 47700
rect 33478 47755 33554 47765
rect 38067 47761 38123 48263
rect 33478 47699 33488 47755
rect 33544 47699 33554 47755
rect 33478 47689 33554 47699
rect 38056 47752 38132 47761
rect 38056 47696 38067 47752
rect 38123 47696 38132 47752
rect 38056 47685 38132 47696
rect 35250 46426 35350 46430
rect 34944 46370 35267 46426
rect 35323 46370 35350 46426
rect 34039 46200 34115 46211
rect 32984 46144 34048 46200
rect 34104 46144 34115 46200
rect 32424 45808 32500 45820
rect 32424 45752 32435 45808
rect 32491 45752 32500 45808
rect 32424 45744 32500 45752
rect 27710 45416 27720 45472
rect 27776 45416 27786 45472
rect 27710 45407 27786 45416
rect 29335 45472 29411 45482
rect 29335 45416 29344 45472
rect 29400 45416 29411 45472
rect 27720 44184 27776 45407
rect 29335 45406 29411 45416
rect 27878 45080 27954 45091
rect 27878 45024 27888 45080
rect 27944 45024 27954 45080
rect 27878 45015 27954 45024
rect 27709 44172 27785 44184
rect 27888 44181 27944 45015
rect 32456 44744 32532 44755
rect 32456 44688 32467 44744
rect 32523 44688 32532 44744
rect 32456 44679 32532 44688
rect 27709 44116 27720 44172
rect 27776 44116 27785 44172
rect 27709 44108 27785 44116
rect 27878 44171 27954 44181
rect 32467 44177 32523 44679
rect 27878 44115 27888 44171
rect 27944 44115 27954 44171
rect 27878 44105 27954 44115
rect 32456 44168 32532 44177
rect 32456 44112 32467 44168
rect 32523 44112 32532 44168
rect 32456 44101 32532 44112
rect 30253 42840 30329 42852
rect 30253 42784 30263 42840
rect 30319 42784 30688 42840
rect 30744 42784 30800 42840
rect 30253 42776 30329 42784
rect 28439 42616 28515 42627
rect 27384 42560 28448 42616
rect 28504 42560 28515 42616
rect 26824 42224 26900 42236
rect 26824 42168 26835 42224
rect 26891 42168 26900 42224
rect 26824 42160 26900 42168
rect 27384 41995 27552 42560
rect 28439 42551 28515 42560
rect 32435 42236 32491 43058
rect 32984 42616 33152 46144
rect 34039 46135 34115 46144
rect 34944 45482 35000 46370
rect 35250 46366 35350 46370
rect 38035 45820 38091 46642
rect 38584 46200 38752 49728
rect 39639 49719 39715 49728
rect 38910 49056 38986 49067
rect 40544 49066 40600 49954
rect 40850 49950 40950 49954
rect 43635 49404 43691 50226
rect 43624 49392 43700 49404
rect 43624 49336 43635 49392
rect 43691 49336 43700 49392
rect 43624 49328 43700 49336
rect 44072 49392 45696 49448
rect 44072 49336 44128 49392
rect 44184 49336 45500 49392
rect 45612 49336 45696 49392
rect 44072 49280 45696 49336
rect 38910 49000 38920 49056
rect 38976 49000 38986 49056
rect 38910 48991 38986 49000
rect 40535 49056 40611 49066
rect 40535 49000 40544 49056
rect 40600 49000 40611 49056
rect 38920 47768 38976 48991
rect 40535 48990 40611 49000
rect 39078 48664 39154 48675
rect 39078 48608 39088 48664
rect 39144 48608 39154 48664
rect 39078 48599 39154 48608
rect 38910 47756 38986 47768
rect 39088 47765 39144 48599
rect 43656 48328 43732 48339
rect 43656 48272 43667 48328
rect 43723 48272 43732 48328
rect 43656 48263 43732 48272
rect 44072 48328 45192 48384
rect 44072 48272 44128 48328
rect 44184 48272 45024 48328
rect 45136 48272 45192 48328
rect 38910 47700 38920 47756
rect 38976 47700 38986 47756
rect 38910 47692 38986 47700
rect 39078 47755 39154 47765
rect 43667 47761 43723 48263
rect 44072 48216 45192 48272
rect 39078 47699 39088 47755
rect 39144 47699 39154 47755
rect 39078 47689 39154 47699
rect 43656 47752 43732 47761
rect 43656 47696 43667 47752
rect 43723 47696 43732 47752
rect 43656 47685 43732 47696
rect 40850 46426 40950 46430
rect 40544 46370 40867 46426
rect 40923 46370 40950 46426
rect 39639 46200 39715 46211
rect 38584 46144 39648 46200
rect 39704 46144 39715 46200
rect 38024 45808 38100 45820
rect 38024 45752 38035 45808
rect 38091 45752 38100 45808
rect 38024 45744 38100 45752
rect 33310 45472 33386 45482
rect 33310 45416 33320 45472
rect 33376 45416 33386 45472
rect 33310 45406 33386 45416
rect 34935 45472 35011 45482
rect 34935 45416 34944 45472
rect 35000 45416 35011 45472
rect 34935 45406 35011 45416
rect 33320 44184 33376 45406
rect 33478 45080 33554 45091
rect 33478 45024 33488 45080
rect 33544 45024 33554 45080
rect 33478 45015 33554 45024
rect 33310 44172 33386 44184
rect 33488 44181 33544 45015
rect 38056 44744 38132 44755
rect 38056 44688 38067 44744
rect 38123 44688 38132 44744
rect 38056 44679 38132 44688
rect 33310 44116 33320 44172
rect 33376 44116 33386 44172
rect 33310 44108 33386 44116
rect 33478 44171 33554 44181
rect 38067 44177 38123 44679
rect 33478 44115 33488 44171
rect 33544 44115 33554 44171
rect 33478 44105 33554 44115
rect 38056 44168 38132 44177
rect 38056 44112 38067 44168
rect 38123 44112 38132 44168
rect 38056 44101 38132 44112
rect 35853 42840 35929 42851
rect 35853 42784 35863 42840
rect 35919 42784 36288 42840
rect 36344 42784 36400 42840
rect 35853 42775 35929 42784
rect 34039 42616 34115 42627
rect 32984 42560 34048 42616
rect 34104 42560 34115 42616
rect 32424 42224 32500 42236
rect 32424 42168 32435 42224
rect 32491 42168 32500 42224
rect 32424 42160 32500 42168
rect 32984 41995 33152 42560
rect 34039 42551 34115 42560
rect 38035 42236 38091 43058
rect 38584 42616 38752 46144
rect 39639 46135 39715 46144
rect 38909 45472 38985 45483
rect 40544 45482 40600 46370
rect 40850 46366 40950 46370
rect 43635 45820 43691 46642
rect 43624 45808 43700 45820
rect 43624 45752 43635 45808
rect 43691 45752 43700 45808
rect 43624 45744 43700 45752
rect 44072 45808 45696 45864
rect 44072 45752 44128 45808
rect 44184 45752 45497 45808
rect 45609 45752 45696 45808
rect 44072 45696 45696 45752
rect 38909 45416 38920 45472
rect 38976 45416 38985 45472
rect 38909 45407 38985 45416
rect 40535 45472 40611 45482
rect 40535 45416 40544 45472
rect 40600 45416 40611 45472
rect 38920 44184 38976 45407
rect 40535 45406 40611 45416
rect 39078 45080 39154 45092
rect 39078 45024 39088 45080
rect 39144 45024 39154 45080
rect 39078 45016 39154 45024
rect 38910 44172 38986 44184
rect 39088 44182 39144 45016
rect 43657 44744 43733 44754
rect 43657 44688 43667 44744
rect 43723 44688 43733 44744
rect 43657 44678 43733 44688
rect 44072 44744 45193 44800
rect 44072 44688 44128 44744
rect 44184 44688 45024 44744
rect 45136 44688 45193 44744
rect 43667 44184 43723 44678
rect 44072 44632 45193 44688
rect 38910 44116 38920 44172
rect 38976 44116 38986 44172
rect 38910 44108 38986 44116
rect 39078 44171 39154 44182
rect 39078 44115 39088 44171
rect 39144 44115 39154 44171
rect 39078 44106 39154 44115
rect 43657 44172 43733 44184
rect 43657 44116 43667 44172
rect 43723 44116 43733 44172
rect 43657 44108 43733 44116
rect 41451 42840 41527 42850
rect 41451 42784 41463 42840
rect 41519 42784 41888 42840
rect 41944 42784 42000 42840
rect 41451 42774 41527 42784
rect 39638 42616 39714 42628
rect 38584 42560 39648 42616
rect 39704 42560 39714 42616
rect 38024 42224 38100 42236
rect 38024 42168 38035 42224
rect 38091 42168 38100 42224
rect 38024 42160 38100 42168
rect 38584 41859 38752 42560
rect 39638 42552 39714 42560
rect 43635 42235 43691 43382
rect 43624 42224 43700 42235
rect 43624 42168 43635 42224
rect 43691 42168 43700 42224
rect 43624 42159 43700 42168
rect 44072 42224 45696 42280
rect 44072 42168 44128 42224
rect 44184 42168 45498 42224
rect 45610 42168 45696 42224
rect 44072 42112 45696 42168
rect 38584 41747 38609 41859
rect 38719 41747 38752 41859
rect 38584 41720 38752 41747
<< via2 >>
rect 2688 42784 2744 42840
rect 8288 42784 8344 42840
rect 13888 42784 13944 42840
rect 19488 42784 19544 42840
rect 25088 42784 25144 42840
rect 30688 42784 30744 42840
rect 36288 42784 36344 42840
rect 41888 42784 41944 42840
rect 38609 41747 38719 41859
<< metal3 >>
rect 38584 41859 38752 41888
rect 38584 41747 38609 41859
rect 38719 41747 38752 41859
rect 38584 41720 38752 41747
<< via3 >>
rect 2632 43232 2744 43344
rect 8232 43232 8344 43344
rect 13832 43232 13944 43344
rect 19432 43232 19544 43344
rect 25032 43232 25144 43344
rect 30632 43232 30744 43344
rect 36232 43232 36344 43344
rect 41832 43232 41944 43344
rect 1232 41776 1344 41888
rect 6832 41776 6944 41888
rect 12432 41776 12544 41888
rect 18032 41776 18144 41888
rect 23632 41776 23744 41888
rect 29232 41776 29344 41888
rect 34832 41776 34944 41888
rect 38609 41747 38719 41859
rect 40432 41776 40544 41888
<< metal4 >>
rect -1792 43344 46256 43456
rect -1792 43232 2632 43344
rect 2744 43232 8232 43344
rect 8344 43232 13832 43344
rect 13944 43232 19432 43344
rect 19544 43232 25032 43344
rect 25144 43232 30632 43344
rect 30744 43232 36232 43344
rect 36344 43232 41832 43344
rect 41944 43232 46256 43344
rect -1792 43120 46256 43232
rect -1792 41888 46256 42000
rect -1792 41776 1232 41888
rect 1344 41776 6832 41888
rect 6944 41776 12432 41888
rect 12544 41776 18032 41888
rect 18144 41776 23632 41888
rect 23744 41776 29232 41888
rect 29344 41776 34832 41888
rect 34944 41859 40432 41888
rect 34944 41776 38609 41859
rect -1792 41747 38609 41776
rect 38719 41776 40432 41859
rect 40544 41776 46256 41888
rect 38719 41747 46256 41776
rect -1792 41664 46256 41747
use unit_cell_aray  unit_cell_array_0
timestamp 1756715696
transform 1 0 5612 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_1
timestamp 1756715696
transform 1 0 11212 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_2
timestamp 1756715696
transform 1 0 16812 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_3
timestamp 1756715696
transform 1 0 22412 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_4
timestamp 1756715696
transform 1 0 28012 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_5
timestamp 1756715696
transform 1 0 33612 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_6
timestamp 1756715696
transform 1 0 39212 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_7
timestamp 1756715696
transform 1 0 12 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_8
timestamp 1756715696
transform 1 0 11212 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_9
timestamp 1756715696
transform 1 0 5612 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_10
timestamp 1756715696
transform 1 0 16812 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_11
timestamp 1756715696
transform 1 0 22412 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_12
timestamp 1756715696
transform 1 0 28012 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_13
timestamp 1756715696
transform 1 0 33612 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_14
timestamp 1756715696
transform 1 0 39212 0 1 42601
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_15
timestamp 1756715696
transform 1 0 12 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_16
timestamp 1756715696
transform 1 0 5612 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_17
timestamp 1756715696
transform 1 0 11212 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_18
timestamp 1756715696
transform 1 0 16812 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_19
timestamp 1756715696
transform 1 0 22412 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_20
timestamp 1756715696
transform 1 0 28012 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_21
timestamp 1756715696
transform 1 0 33612 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_22
timestamp 1756715696
transform 1 0 39212 0 1 49769
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_23
timestamp 1756715696
transform 1 0 12 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_24
timestamp 1756715696
transform 1 0 5612 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_25
timestamp 1756715696
transform 1 0 11212 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_26
timestamp 1756715696
transform 1 0 16812 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_27
timestamp 1756715696
transform 1 0 22412 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_28
timestamp 1756715696
transform 1 0 28012 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_29
timestamp 1756715696
transform 1 0 33612 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_30
timestamp 1756715696
transform 1 0 39212 0 1 53353
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_31
timestamp 1756715696
transform 1 0 12 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_32
timestamp 1756715696
transform 1 0 11212 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_33
timestamp 1756715696
transform 1 0 5612 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_34
timestamp 1756715696
transform 1 0 16812 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_35
timestamp 1756715696
transform 1 0 22412 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_36
timestamp 1756715696
transform 1 0 33612 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_37
timestamp 1756715696
transform 1 0 28012 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_38
timestamp 1756715696
transform 1 0 39212 0 1 56937
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_39
timestamp 1756715696
transform 1 0 12 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_40
timestamp 1756715696
transform 1 0 12 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_41
timestamp 1756715696
transform 1 0 12 0 1 46185
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_42
timestamp 1756715696
transform 1 0 5612 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_43
timestamp 1756715696
transform 1 0 11212 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_44
timestamp 1756715696
transform 1 0 11212 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_45
timestamp 1756715696
transform 1 0 5612 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_46
timestamp 1756715696
transform 1 0 16812 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_47
timestamp 1756715696
transform 1 0 16812 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_48
timestamp 1756715696
transform 1 0 22412 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_49
timestamp 1756715696
transform 1 0 22412 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_50
timestamp 1756715696
transform 1 0 28012 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_51
timestamp 1756715696
transform 1 0 33612 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_52
timestamp 1756715696
transform 1 0 33612 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_53
timestamp 1756715696
transform 1 0 28012 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_54
timestamp 1756715696
transform 1 0 39212 0 1 64105
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_55
timestamp 1756715696
transform 1 0 39212 0 1 60521
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_56
timestamp 1756715696
transform 1 0 12 0 1 67689
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_57
timestamp 1756715696
transform 1 0 5612 0 1 67689
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_58
timestamp 1756715696
transform 1 0 11212 0 1 67689
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_59
timestamp 1756715696
transform 1 0 16812 0 1 67689
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_60
timestamp 1756715696
transform 1 0 22412 0 1 67689
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_61
timestamp 1756715696
transform 1 0 28012 0 1 67689
box -12 -1288 4835 2603
use unit_cell_aray  unit_cell_array_62
timestamp 1756715696
transform 1 0 33612 0 1 67689
box -12 -1288 4835 2603
<< labels >>
flabel metal1 44408 41776 44744 70565 1 FreeSans 8000 0 0 0 OUTP
port 16 n
flabel space 44912 69219 45248 70567 1 FreeSans 8000 0 0 0 OUTN
port 17 n
rlabel metal1 44912 41776 45248 70565 1 OUTN
port 17 n
flabel metal1 -168 45360 1344 45528 1 FreeSans 3200 0 0 0 D1
port 1 n
flabel metal1 -224 48944 1344 49112 1 FreeSans 3200 0 0 0 D2
port 2 n
flabel metal1 -224 52528 1344 52696 1 FreeSans 3200 0 0 0 D3
port 3 n
flabel metal1 -224 56112 1344 56280 1 FreeSans 3200 0 0 0 D4
port 4 n
flabel metal1 -224 59696 1344 59864 1 FreeSans 3200 0 0 0 D5
port 5 n
flabel metal1 -224 63280 1344 63448 1 FreeSans 3200 0 0 0 D6
port 6 n
flabel metal1 -224 66864 1344 67032 1 FreeSans 3200 0 0 0 D7
port 7 n
flabel metal2 -616 69561 -448 70461 1 FreeSans 3200 0 0 0 C1
port 8 n
flabel metal2 4984 69499 5152 70399 1 FreeSans 3200 0 0 0 C2
port 9 n
flabel metal2 10584 69609 10752 70509 1 FreeSans 3200 0 0 0 C3
port 10 n
flabel metal2 21784 69438 21952 70338 1 FreeSans 3200 0 0 0 C5
port 12 n
flabel metal2 27384 69435 27552 70335 1 FreeSans 3200 0 0 0 C6
port 13 n
flabel metal2 32984 69565 33152 70465 1 FreeSans 3200 0 0 0 C7
port 14 n
flabel metal1 -952 41776 -784 70461 1 FreeSans 3200 0 0 0 CLK
port 15 n
flabel metal1 45416 41776 45752 70565 1 FreeSans 3200 0 0 0 VBIAS
port 18 n
flabel metal2 16184 69357 16352 70265 1 FreeSans 3200 0 0 0 C4
port 11 n
flabel metal4 -1792 43120 46256 43456 1 FreeSans 8000 0 0 0 VDD
port 19 n
flabel metal4 -1792 41664 46256 42000 1 FreeSans 8000 0 0 0 VSS
port 20 n
<< end >>
