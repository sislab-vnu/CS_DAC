VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CS_Switch_1x
  CLASS BLOCK ;
  FOREIGN CS_Switch_1x ;
  ORIGIN 1.630 9.445 ;
  SIZE 8.565 BY 4.325 ;
  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.061600 ;
    PORT
      LAYER Metal1 ;
        RECT -0.260 -7.100 -0.030 -6.450 ;
    END
  END INP
  PIN INN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.061600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.890 -7.100 1.120 -6.450 ;
    END
  END INN
  PIN OUTP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT -0.845 -7.250 -0.555 -6.225 ;
        RECT -0.895 -7.635 -0.515 -7.250 ;
    END
  END OUTP
  PIN OUTN
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.425 -7.265 1.715 -6.225 ;
        RECT 1.375 -7.650 1.755 -7.265 ;
    END
  END OUTN
  PIN VBIAS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.710 -7.230 5.640 -6.875 ;
    END
  END VBIAS
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.965 -7.620 6.345 -7.235 ;
        RECT 6.005 -8.450 6.310 -7.620 ;
        RECT -1.145 -9.025 6.415 -8.450 ;
        RECT -1.145 -9.030 0.380 -9.025 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -1.630 -9.445 6.935 -5.120 ;
    END
  END VPW
  OBS
      LAYER Metal1 ;
        RECT 0.240 -7.635 0.620 -7.250 ;
        RECT 2.170 -7.620 2.550 -7.235 ;
        RECT 0.280 -7.935 0.570 -7.635 ;
        RECT 2.235 -7.935 2.525 -7.620 ;
        RECT 0.280 -8.170 2.525 -7.935 ;
  END
END CS_Switch_1x
END LIBRARY

