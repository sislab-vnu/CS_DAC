VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CS_Switch_16x
  CLASS BLOCK ;
  FOREIGN CS_Switch_16x ;
  ORIGIN -5.110 2.435 ;
  SIZE 5.170 BY 3.765 ;
  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 -0.655 6.280 -0.620 ;
        RECT 5.425 -0.985 6.280 -0.655 ;
        RECT 5.900 -1.000 6.280 -0.985 ;
    END
  END INP
  PIN INN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 0.520 6.280 0.540 ;
        RECT 5.425 0.190 6.280 0.520 ;
        RECT 5.900 0.160 6.280 0.190 ;
    END
  END INN
  PIN OUTP
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.234000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.630 -1.080 7.010 -1.040 ;
        RECT 6.520 -1.390 7.280 -1.080 ;
        RECT 6.630 -1.420 7.010 -1.390 ;
    END
  END OUTP
  PIN OUTN
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.630 0.930 7.010 0.960 ;
        RECT 6.510 0.620 7.310 0.930 ;
        RECT 6.630 0.580 7.010 0.620 ;
    END
  END OUTN
  PIN VBIAS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.260 1.015 8.640 1.050 ;
        RECT 8.040 0.685 8.845 1.015 ;
        RECT 8.260 0.670 8.640 0.685 ;
    END
  END VBIAS
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 -0.420 9.480 -0.040 ;
        RECT 9.170 -1.660 9.410 -0.420 ;
        RECT 5.880 -2.185 9.830 -1.660 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 5.110 0.930 10.280 1.330 ;
        RECT 5.110 0.620 6.510 0.930 ;
        RECT 6.620 0.730 7.020 0.930 ;
        RECT 6.520 0.620 7.120 0.730 ;
        RECT 7.310 0.620 10.280 0.930 ;
        RECT 5.110 -1.075 10.280 0.620 ;
        RECT 5.110 -1.190 7.120 -1.075 ;
        RECT 5.110 -1.390 6.520 -1.190 ;
        RECT 6.620 -1.390 7.020 -1.190 ;
        RECT 7.320 -1.390 10.280 -1.075 ;
        RECT 5.110 -2.435 10.280 -1.390 ;
    END
  END VPW
  OBS
      LAYER Metal1 ;
        RECT 6.630 -0.110 7.010 -0.040 ;
        RECT 7.410 -0.110 7.790 -0.040 ;
        RECT 6.630 -0.350 7.790 -0.110 ;
        RECT 6.630 -0.420 7.010 -0.350 ;
        RECT 7.410 -0.420 7.790 -0.350 ;
  END
END CS_Switch_16x
END LIBRARY

