* NGSPICE file created from CS_Switch_1x1.ext - technology: gf180mcuD

.subckt CS_Switch_1x1 INP INN OUTP OUTN VBIAS VSS
X0 a_668_n40# VSS.t11 a_440_n224# VSS.t10 nfet_03v3 ad=50.6f pd=0.9u as=0.1452p ps=1.465u w=0.22u l=0.28u
X1 a_668_n224# VSS.t9 a_440_n224# VSS.t10 nfet_03v3 ad=50.6f pd=0.9u as=0.1452p ps=1.465u w=0.22u l=0.28u
X2 a_440_n224# VBIAS.t0 a_56_n40# VSS.t0 nfet_03v3 ad=0.1452p pd=1.465u as=0.1516p ps=1.64u w=0.22u l=0.28u
X3 VSS.t8 VSS.t7 a_n228_n224# VSS.t6 nfet_03v3 ad=94.5f pd=0.99u as=50.6f ps=0.9u w=0.22u l=0.28u
X4 OUTN.t0 INN.t0 a_56_n40# VSS.t3 nfet_03v3 ad=0.182p pd=1.8u as=86.8f ps=0.92u w=0.22u l=0.28u
X5 a_440_n224# VBIAS.t1 VSS.t2 VSS.t1 nfet_03v3 ad=0.1452p pd=1.465u as=94.5f ps=0.99u w=0.22u l=2.2u
X6 a_56_n40# INP.t0 OUTP.t0 VSS.t4 nfet_03v3 ad=86.8f pd=0.92u as=0.1053p ps=1.03u w=0.22u l=0.28u
X7 OUTP.t1 VSS.t5 a_n228_n40# VSS.t6 nfet_03v3 ad=0.1053p pd=1.03u as=50.6f ps=0.9u w=0.22u l=0.28u
R0 VSS VSS.t1 1253.86
R1 VSS.t4 VSS.t6 912.809
R2 VSS.t3 VSS.t4 842.593
R3 VSS.n1 VSS 371.142
R4 VSS VSS.t10 235.726
R5 VSS.t0 VSS 150.464
R6 VSS.t1 VSS.t3 120.371
R7 VSS.n1 VSS.t0 95.2937
R8 VSS.t9 VSS.t11 23.9862
R9 VSS.t7 VSS.t5 23.9862
R10 VSS.n2 VSS.t9 20.5166
R11 VSS.n3 VSS.t7 20.4235
R12 VSS.n2 VSS.n1 10.4005
R13 VSS.n0 VSS.t8 8.01868
R14 VSS VSS.n0 6.40615
R15 VSS.n0 VSS.t2 6.01414
R16 VSS VSS.n2 0.439059
R17 VSS VSS.n3 0.0744831
R18 VSS.n3 VSS 0.0378729
R19 VBIAS.t0 VBIAS.t1 43.9669
R20 VBIAS VBIAS.t0 22.6455
R21 INN INN.t0 22.6455
R22 OUTN.n0 OUTN.t0 12.3141
R23 OUTN OUTN.n0 0.0455
R24 OUTN.n0 OUTN 0.0455
R25 INP INP.t0 22.6455
R26 OUTP.n0 OUTP.t1 6.87323
R27 OUTP OUTP.n0 6.3455
R28 OUTP.n0 OUTP.t0 6.01414
C0 a_668_n224# VSS 8.29e-19
C1 OUTP a_n228_n40# 7.7e-19
C2 OUTP OUTN 6.32e-19
C3 OUTP INN 7.62e-20
C4 OUTP VSS 0.02973f
C5 OUTN VBIAS 0.001717f
C6 OUTN a_56_n40# 0.164087f
C7 OUTN INP 7.62e-20
C8 VBIAS a_440_n224# 0.001013f
C9 a_56_n40# a_440_n224# 0.00171f
C10 INN VBIAS 0.041164f
C11 INN a_56_n40# 0.029406f
C12 VBIAS VSS 0.580307f
C13 INN INP 0.060872f
C14 a_56_n40# VSS 0.150521f
C15 VSS INP 0.132936f
C16 a_n228_n40# VSS 2.43e-19
C17 a_n228_n224# VSS 3.61e-19
C18 OUTN INN 0.003858f
C19 OUTP a_56_n40# 0.029701f
C20 OUTN VSS 4.68e-20
C21 OUTP INP 0.003858f
C22 a_440_n224# VSS 0.006325f
C23 INN VSS 0.113785f
C24 VBIAS a_56_n40# 0.047893f
C25 VBIAS INP 0.019271f
C26 a_56_n40# INP 0.003069f
C27 a_668_n40# VSS 5.59e-19
C28 OUTN VSUBS 0.018808f
C29 OUTP VSUBS 0.030912f
C30 VBIAS VSUBS 0.358538f
C31 INN VSUBS 0.064325f
C32 INP VSUBS 0.079541f
C33 VSS VSUBS 0.5802f
C34 a_56_n40# VSUBS 0.105866f
.ends

