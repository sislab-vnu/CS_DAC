magic
tech gf180mcuD
magscale 1 10
timestamp 1755157607
<< pwell >>
rect 3920 -591 5359 -73
rect 3920 -1029 6677 -591
rect 8245 -701 8592 -591
rect 8673 -701 9552 -591
rect 8245 -1029 9552 -701
rect 3920 -1547 5359 -1029
rect 3920 -1985 6677 -1547
rect 8245 -1662 8584 -1547
rect 8700 -1662 9566 -1547
rect 8245 -1985 9566 -1662
rect 3920 -2511 5359 -1985
rect 3920 -2963 5535 -2511
rect 3920 -3482 5359 -2963
rect 3920 -3920 6677 -3482
rect 8245 -3621 8553 -3482
rect 8720 -3621 9668 -3482
rect 8245 -3920 9668 -3621
rect 3920 -3993 5359 -3920
<< metal1 >>
rect 2352 -348 2688 56
rect 2914 -301 2968 -237
rect 3080 -301 5062 -237
rect 4998 -302 5062 -301
rect 2352 -412 4651 -348
rect 2352 -1273 2688 -412
rect 4589 -682 4651 -412
rect 4998 -609 5063 -302
rect 4972 -674 5063 -609
rect 5983 -602 6312 -519
rect 9800 -513 10080 -280
rect 9441 -589 10080 -513
rect 5135 -883 5275 -881
rect 5135 -1001 5447 -883
rect 2874 -1224 2968 -1160
rect 3081 -1224 5037 -1160
rect 2352 -1337 4626 -1273
rect 2352 -2225 2688 -1337
rect 4563 -1599 4626 -1337
rect 4975 -1362 5037 -1224
rect 4974 -1599 5037 -1362
rect 5989 -1558 6309 -1475
rect 9800 -1469 10080 -589
rect 9457 -1546 10080 -1469
rect 5157 -1959 5446 -1839
rect 5237 -1960 5319 -1959
rect 2900 -2178 2968 -2116
rect 3080 -2178 4780 -2116
rect 2900 -2179 4780 -2178
rect 4719 -2212 4780 -2179
rect 2352 -2289 4374 -2225
rect 2352 -3317 2688 -2289
rect 4311 -2554 4374 -2289
rect 4719 -2554 4782 -2287
rect 5986 -2521 6326 -2438
rect 9800 -2432 10080 -1546
rect 9456 -2508 10080 -2432
rect 5154 -2922 5498 -2802
rect 2897 -3148 2968 -3083
rect 3080 -3148 5173 -3083
rect 2352 -3382 4706 -3317
rect 2352 -4032 2688 -3382
rect 4301 -3434 4464 -3431
rect 4301 -3487 4326 -3434
rect 4451 -3487 4464 -3434
rect 4301 -3495 4464 -3487
rect 4641 -3626 4706 -3382
rect 5108 -3623 5173 -3148
rect 5989 -3493 6327 -3410
rect 9800 -3404 10080 -2508
rect 9456 -3480 10080 -3404
rect 9800 -3640 10080 -3480
rect 5232 -3894 5451 -3774
<< via1 >>
rect 2968 -301 3080 -237
rect 4407 -548 4463 -496
rect 4711 -547 4765 -494
rect 4878 -548 4936 -494
rect 6341 -460 6481 -374
rect 5581 -634 5641 -547
rect 8600 -685 8663 -446
rect 2968 -1224 3081 -1160
rect 4384 -1464 4437 -1412
rect 4686 -1466 4741 -1413
rect 4863 -1467 4917 -1413
rect 6351 -1406 6474 -1340
rect 5581 -1590 5641 -1505
rect 8609 -1638 8666 -1385
rect 2968 -2178 3080 -2116
rect 4127 -2420 4181 -2368
rect 4429 -2421 4484 -2367
rect 4606 -2421 4661 -2367
rect 4911 -2420 4965 -2367
rect 6357 -2371 6473 -2302
rect 5582 -2554 5642 -2470
rect 8609 -2600 8665 -2346
rect 2968 -3148 3080 -3083
rect 4326 -3487 4451 -3434
rect 4767 -3505 4823 -3449
rect 4994 -3506 5052 -3448
rect 6361 -3341 6475 -3281
rect 5582 -3525 5642 -3445
rect 8607 -3577 8665 -3324
<< metal2 >>
rect 2856 -237 3192 56
rect 2856 -301 2968 -237
rect 3080 -301 3192 -237
rect 2856 -1160 3192 -301
rect 4701 -355 5457 -354
rect 6305 -355 6521 -348
rect 4701 -374 6521 -355
rect 4701 -423 6341 -374
rect 4701 -481 4780 -423
rect 5001 -424 6341 -423
rect 6305 -460 6341 -424
rect 6481 -460 6521 -374
rect 6305 -477 6521 -460
rect 8592 -446 8673 -401
rect 4395 -484 4475 -481
rect 3404 -559 3462 -484
rect 3580 -496 4475 -484
rect 3580 -548 4407 -496
rect 4463 -548 4475 -496
rect 3580 -559 4475 -548
rect 4395 -561 4475 -559
rect 4699 -494 4780 -481
rect 4699 -547 4711 -494
rect 4765 -508 4780 -494
rect 4867 -490 4947 -481
rect 4867 -494 5662 -490
rect 4765 -547 4779 -508
rect 4699 -561 4779 -547
rect 4867 -548 4878 -494
rect 4936 -547 5662 -494
rect 4936 -548 5581 -547
rect 4867 -559 5581 -548
rect 4867 -561 4947 -559
rect 5551 -634 5581 -559
rect 5641 -559 5662 -547
rect 5641 -634 5661 -559
rect 5551 -648 5661 -634
rect 8592 -685 8600 -446
rect 8663 -685 8673 -446
rect 8592 -701 8673 -685
rect 2856 -1224 2968 -1160
rect 3081 -1224 3192 -1160
rect 2856 -2116 3192 -1224
rect 4675 -1340 6524 -1271
rect 4675 -1341 6351 -1340
rect 4675 -1399 4751 -1341
rect 4370 -1402 4450 -1399
rect 3410 -1403 4450 -1402
rect 3410 -1477 3472 -1403
rect 3584 -1412 4450 -1403
rect 3584 -1464 4384 -1412
rect 4437 -1464 4450 -1412
rect 3584 -1477 4450 -1464
rect 4370 -1479 4450 -1477
rect 4674 -1413 4754 -1399
rect 4674 -1466 4686 -1413
rect 4741 -1466 4754 -1413
rect 4674 -1479 4754 -1466
rect 4850 -1409 4930 -1399
rect 6307 -1406 6351 -1341
rect 6474 -1341 6524 -1340
rect 6474 -1406 6523 -1341
rect 4850 -1413 5663 -1409
rect 4850 -1467 4863 -1413
rect 4917 -1467 5663 -1413
rect 6307 -1433 6523 -1406
rect 8594 -1385 8675 -1357
rect 4850 -1479 5663 -1467
rect 5555 -1505 5663 -1479
rect 5555 -1590 5581 -1505
rect 5641 -1590 5663 -1505
rect 5555 -1604 5663 -1590
rect 8594 -1638 8609 -1385
rect 8666 -1638 8675 -1385
rect 8594 -1657 8675 -1638
rect 2856 -2178 2968 -2116
rect 3080 -2178 3192 -2116
rect 2856 -3083 3192 -2178
rect 4419 -2159 6523 -2089
rect 4419 -2354 4486 -2159
rect 4596 -2290 5640 -2220
rect 4596 -2354 4672 -2290
rect 4116 -2366 4192 -2356
rect 3446 -2432 3472 -2366
rect 3583 -2368 4192 -2366
rect 3583 -2420 4127 -2368
rect 4181 -2420 4192 -2368
rect 3583 -2432 4192 -2420
rect 4418 -2367 4498 -2354
rect 4418 -2421 4429 -2367
rect 4484 -2421 4498 -2367
rect 4119 -2693 4188 -2432
rect 4418 -2434 4498 -2421
rect 4594 -2367 4674 -2354
rect 4594 -2421 4606 -2367
rect 4661 -2421 4674 -2367
rect 4594 -2434 4674 -2421
rect 4898 -2367 4978 -2354
rect 4898 -2420 4911 -2367
rect 4965 -2420 4978 -2367
rect 4898 -2434 4978 -2420
rect 4904 -2693 4973 -2434
rect 5555 -2449 5640 -2290
rect 6308 -2267 6523 -2159
rect 6308 -2302 6524 -2267
rect 6308 -2371 6357 -2302
rect 6473 -2371 6524 -2302
rect 6308 -2396 6524 -2371
rect 8595 -2346 8676 -2320
rect 5555 -2470 5669 -2449
rect 5555 -2554 5582 -2470
rect 5642 -2554 5669 -2470
rect 5555 -2567 5669 -2554
rect 5555 -2568 5666 -2567
rect 8595 -2600 8609 -2346
rect 8665 -2600 8676 -2346
rect 8595 -2620 8676 -2600
rect 4119 -2762 4973 -2693
rect 2856 -3148 2968 -3083
rect 3080 -3148 3192 -3083
rect 2856 -4032 3192 -3148
rect 4757 -3281 6524 -3219
rect 4757 -3289 6361 -3281
rect 3398 -3496 3433 -3430
rect 3589 -3434 4465 -3430
rect 3589 -3487 4326 -3434
rect 4451 -3487 4465 -3434
rect 4757 -3437 4827 -3289
rect 6308 -3341 6361 -3289
rect 6475 -3341 6524 -3281
rect 6308 -3368 6524 -3341
rect 8595 -3324 8676 -3292
rect 3589 -3496 4465 -3487
rect 4755 -3449 4835 -3437
rect 4755 -3505 4767 -3449
rect 4823 -3505 4835 -3449
rect 4755 -3517 4835 -3505
rect 4983 -3445 5063 -3437
rect 5563 -3445 5664 -3429
rect 4983 -3448 5582 -3445
rect 4983 -3506 4994 -3448
rect 5052 -3506 5582 -3448
rect 4983 -3515 5582 -3506
rect 4983 -3517 5063 -3515
rect 5563 -3525 5582 -3515
rect 5642 -3525 5664 -3445
rect 5563 -3539 5664 -3525
rect 8595 -3577 8607 -3324
rect 8665 -3577 8676 -3324
rect 8595 -3592 8676 -3577
<< via2 >>
rect 3462 -559 3580 -484
rect 3472 -1477 3584 -1403
rect 3472 -2432 3583 -2366
rect 3433 -3496 3589 -3430
<< metal3 >>
rect 3360 -484 3696 56
rect 3360 -559 3462 -484
rect 3580 -559 3696 -484
rect 3360 -1403 3696 -559
rect 3360 -1477 3472 -1403
rect 3584 -1477 3696 -1403
rect 3360 -2366 3696 -1477
rect 3360 -2432 3472 -2366
rect 3583 -2432 3696 -2366
rect 3360 -3430 3696 -2432
rect 3360 -3496 3433 -3430
rect 3589 -3496 3696 -3430
rect 3360 -4032 3696 -3496
use CS_Switch_1x1  CS_Switch_1x1_0
timestamp 1754893325
transform -1 0 4935 0 1 -627
box -306 -434 837 214
use CS_Switch_2x2  CS_Switch_2x2_0
timestamp 1754896527
transform -1 0 4894 0 1 -1563
box -356 -436 795 224
use CS_Switch_4x2  CS_Switch_4x2_0
timestamp 1754896551
transform 1 0 4140 0 1 -2778
box -304 -185 1117 488
use CS_Switch_8x2  CS_Switch_8x2_0
timestamp 1754903761
transform -1 0 5779 0 1 -5007
box 426 1024 1804 1719
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform -1 0 9590 0 1 -2862
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_1
timestamp 1753044640
transform -1 0 9587 0 1 -943
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_2
timestamp 1753044640
transform -1 0 9589 0 1 -1899
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  gf180mcu_fd_sc_mcu7t5v0__dffq_2_3
timestamp 1753044640
transform -1 0 9590 0 1 -3834
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform -1 0 6118 0 1 -2862
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_1
timestamp 1753044640
transform -1 0 6117 0 1 -943
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_2
timestamp 1753044640
transform -1 0 6117 0 1 -1899
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_3
timestamp 1753044640
transform -1 0 6118 0 1 -3834
box -86 -86 758 870
<< labels >>
flabel metal2 8592 -701 8673 -401 1 FreeSans 400 0 0 0 D1
port 1 n
flabel metal2 8594 -1657 8675 -1357 1 FreeSans 400 0 0 0 D2
port 2 n
flabel metal2 8595 -2620 8676 -2320 1 FreeSans 400 0 0 0 D3
port 3 n
flabel metal2 8595 -3592 8676 -3292 1 FreeSans 400 0 0 0 D4
port 4 n
<< end >>
