magic
tech gf180mcuD
magscale 1 10
timestamp 1755162181
<< nwell >>
rect 18259 -970 18308 -918
rect 3478 -6067 3590 -5601
rect 4037 -5666 4089 -5614
rect 2863 -11970 2929 -11959
rect 37953 -14068 38013 -14012
<< pwell >>
rect 3478 -5601 3590 -5163
<< mvpmos >>
rect 2863 -11970 2929 -11959
<< polysilicon >>
rect 4037 -5666 4089 -5614
rect 37953 -14068 38013 -14012
<< metal1 >>
rect 2800 2497 32984 2632
rect 2800 2494 28000 2497
rect 2800 2492 13496 2494
rect 2800 2436 3696 2492
rect 3752 2436 8568 2492
rect 8624 2438 13496 2492
rect 13552 2492 28000 2494
rect 13552 2491 23184 2492
rect 13552 2438 18256 2491
rect 8624 2436 18256 2438
rect 2800 2435 18256 2436
rect 18312 2436 23184 2491
rect 23240 2441 28000 2492
rect 28056 2464 32984 2497
rect 28056 2441 32872 2464
rect 23240 2436 32872 2441
rect 18312 2435 32872 2436
rect 2800 2408 32872 2435
rect 32928 2408 32984 2464
rect 2800 2296 32984 2408
rect 11997 1323 12498 1400
rect 13020 1361 13787 1438
rect 3483 1195 6151 1315
rect 13710 1273 13787 1361
rect 17975 1343 18634 1421
rect 21615 1383 22231 1457
rect 22722 1387 23474 1461
rect 13710 1206 13719 1273
rect 13776 1206 13787 1273
rect 13710 1181 13787 1206
rect 18556 1254 18634 1343
rect 18556 1188 18565 1254
rect 18626 1188 18634 1254
rect 23399 1298 23474 1387
rect 27799 1334 28354 1417
rect 31308 1380 31922 1470
rect 32432 1350 33173 1440
rect 23399 1229 23407 1298
rect 23464 1229 23474 1298
rect 23399 1192 23474 1229
rect 28268 1287 28354 1334
rect 28268 1224 28280 1287
rect 28337 1224 28354 1287
rect 28268 1196 28354 1224
rect 33082 1262 33173 1350
rect 33082 1202 33095 1262
rect 33156 1202 33173 1262
rect 18556 1166 18634 1188
rect 33082 1179 33173 1202
rect 3099 805 4095 870
rect 4028 537 4095 805
rect 43568 672 43904 1400
rect 4028 485 4032 537
rect 4088 485 4095 537
rect 8008 504 43904 672
rect 4028 472 4095 485
rect 3487 291 3714 411
rect 4812 84 5370 103
rect 4437 80 5370 84
rect 4406 39 5370 80
rect 4406 37 4852 39
rect 4406 16 4437 37
rect 4929 -73 5485 -9
rect 3494 -613 3805 -373
rect 4929 -576 4993 -73
rect 3681 -983 3700 -907
rect 3768 -983 3807 -907
rect 8040 -965 8116 504
rect 9658 91 10300 103
rect 9283 82 10300 91
rect 9212 39 10300 82
rect 9212 37 9698 39
rect 9212 18 9283 37
rect 9775 -73 10705 -9
rect 8872 -280 8944 -127
rect 9775 -387 9839 -73
rect 8559 -983 8574 -907
rect 8632 -983 8738 -907
rect 12886 -965 12962 504
rect 14504 91 15146 103
rect 14058 39 15146 91
rect 14058 37 14544 39
rect 14058 27 14129 37
rect 14621 -73 15551 -9
rect 13718 -188 13790 -152
rect 14621 -613 14685 -73
rect 17732 -965 17808 504
rect 19350 90 19992 103
rect 18904 39 19992 90
rect 18904 37 19390 39
rect 18904 26 18975 37
rect 19467 -73 20397 -9
rect 19467 -613 19531 -73
rect 18247 -918 18359 -907
rect 18247 -970 18259 -918
rect 18311 -970 18359 -918
rect 22578 -965 22654 504
rect 24196 94 24838 103
rect 23750 39 24838 94
rect 23750 37 24236 39
rect 23750 30 23821 37
rect 24313 -73 25243 -9
rect 24313 -613 24377 -73
rect 27424 -965 27500 504
rect 29042 93 29684 103
rect 28596 39 29684 93
rect 28596 37 29082 39
rect 28596 29 28667 37
rect 29159 -73 30089 -9
rect 29159 -613 29223 -73
rect 27978 -918 28083 -907
rect 18247 -983 18359 -970
rect 27978 -971 28001 -918
rect 28056 -971 28083 -918
rect 32270 -965 32346 504
rect 33888 93 34530 103
rect 33442 39 34530 93
rect 33442 37 33928 39
rect 33442 29 33513 37
rect 34005 -73 34935 -9
rect 33102 -183 33174 -153
rect 34005 -613 34069 -73
rect 32849 -915 32941 -907
rect 27978 -983 28083 -971
rect 32849 -972 32869 -915
rect 32932 -972 32941 -915
rect 37116 -965 37192 504
rect 37746 148 37796 340
rect 38734 95 39376 103
rect 38287 39 39376 95
rect 38287 37 38773 39
rect 38287 31 38359 37
rect 38851 -73 39781 -9
rect 38851 -613 38915 -73
rect 41962 -965 42038 504
rect 32849 -983 32941 -972
rect 3511 -1397 3753 -1277
rect 43568 -2128 43904 504
rect 8008 -2296 43904 -2128
rect 4846 -2702 5484 -2697
rect 4846 -2755 4893 -2702
rect 4956 -2755 5484 -2702
rect 4846 -2761 5484 -2755
rect 4406 -2873 5280 -2809
rect 3497 -3413 3749 -3293
rect 3671 -3783 3687 -3707
rect 3755 -3783 3835 -3707
rect 8040 -3765 8116 -2296
rect 9713 -2701 10374 -2697
rect 9713 -2754 9772 -2701
rect 9834 -2754 10374 -2701
rect 9713 -2761 10374 -2754
rect 9230 -2873 10144 -2809
rect 8549 -3783 8568 -3707
rect 8628 -3783 8728 -3707
rect 12886 -3765 12962 -2296
rect 14549 -2705 15056 -2697
rect 14549 -2757 14580 -2705
rect 14645 -2757 15056 -2705
rect 14549 -2761 15056 -2757
rect 14093 -2873 15025 -2809
rect 17732 -3765 17808 -2296
rect 19371 -2706 19899 -2697
rect 19371 -2758 19458 -2706
rect 19521 -2758 19899 -2706
rect 19371 -2761 19899 -2758
rect 18905 -2873 20398 -2809
rect 18248 -3719 18368 -3707
rect 18248 -3773 18261 -3719
rect 18319 -3773 18368 -3719
rect 22578 -3765 22654 -2296
rect 24212 -2703 24784 -2697
rect 24212 -2756 24269 -2703
rect 24334 -2756 24784 -2703
rect 24212 -2761 24784 -2756
rect 23789 -2873 25283 -2809
rect 18248 -3783 18368 -3773
rect 27424 -3765 27500 -2296
rect 29050 -2705 29560 -2697
rect 29050 -2758 29145 -2705
rect 29206 -2758 29560 -2705
rect 29050 -2761 29560 -2758
rect 28617 -2873 30052 -2809
rect 27980 -3718 28079 -3707
rect 27980 -3770 27993 -3718
rect 28049 -3770 28079 -3718
rect 32270 -3765 32346 -2296
rect 33926 -2705 34786 -2697
rect 33926 -2757 33989 -2705
rect 34051 -2757 34786 -2705
rect 33926 -2761 34786 -2757
rect 33465 -2873 34789 -2809
rect 32854 -3714 32935 -3707
rect 27980 -3783 28079 -3770
rect 32854 -3774 32869 -3714
rect 32932 -3774 32935 -3714
rect 37116 -3765 37192 -2296
rect 38769 -2706 39440 -2697
rect 38769 -2758 38833 -2706
rect 38894 -2758 39440 -2706
rect 38769 -2761 39440 -2758
rect 38350 -2873 39689 -2809
rect 41962 -3765 42038 -2296
rect 32854 -3783 32935 -3774
rect 3468 -4197 3720 -4077
rect 43568 -4928 43904 -2296
rect 8008 -5096 43904 -4928
rect 3370 -5309 3709 -5189
rect 4846 -5502 5484 -5497
rect 4846 -5555 4893 -5502
rect 4956 -5555 5484 -5502
rect 4846 -5561 5484 -5555
rect 4406 -5673 5280 -5609
rect 3294 -6213 3701 -5973
rect 3678 -6583 3691 -6507
rect 3750 -6583 3829 -6507
rect 8040 -6565 8116 -5096
rect 9713 -5501 10374 -5497
rect 9713 -5554 9772 -5501
rect 9834 -5554 10374 -5501
rect 9713 -5561 10374 -5554
rect 9230 -5673 10144 -5609
rect 8548 -6583 8565 -6507
rect 8624 -6583 8714 -6507
rect 12886 -6565 12962 -5096
rect 14549 -5505 15056 -5497
rect 14549 -5557 14580 -5505
rect 14645 -5557 15056 -5505
rect 14549 -5561 15056 -5557
rect 14093 -5673 15025 -5609
rect 17732 -6565 17808 -5096
rect 19371 -5506 19899 -5497
rect 19371 -5558 19458 -5506
rect 19521 -5558 19899 -5506
rect 19371 -5561 19899 -5558
rect 18905 -5673 20398 -5609
rect 18246 -6520 18369 -6507
rect 18246 -6573 18257 -6520
rect 18315 -6573 18369 -6520
rect 22578 -6565 22654 -5096
rect 24212 -5503 24784 -5497
rect 24212 -5556 24269 -5503
rect 24334 -5556 24784 -5503
rect 24212 -5561 24784 -5556
rect 23789 -5673 25283 -5609
rect 27424 -6565 27500 -5096
rect 29050 -5505 29560 -5497
rect 29050 -5558 29145 -5505
rect 29206 -5558 29560 -5505
rect 29050 -5561 29560 -5558
rect 28617 -5673 30052 -5609
rect 27973 -6519 28070 -6507
rect 18246 -6583 18369 -6573
rect 27973 -6574 27989 -6519
rect 28042 -6574 28070 -6519
rect 32270 -6565 32346 -5096
rect 33926 -5505 34767 -5497
rect 33926 -5557 33989 -5505
rect 34051 -5557 34767 -5505
rect 33926 -5561 34767 -5557
rect 33465 -5673 34789 -5609
rect 32858 -6518 32939 -6507
rect 27973 -6583 28070 -6574
rect 32858 -6573 32870 -6518
rect 32933 -6573 32939 -6518
rect 37116 -6565 37192 -5096
rect 37745 -5452 37796 -5284
rect 38769 -5506 39440 -5497
rect 38769 -5558 38833 -5506
rect 38894 -5558 39440 -5506
rect 38769 -5561 39440 -5558
rect 38350 -5673 39689 -5609
rect 41962 -6565 42038 -5096
rect 32858 -6583 32939 -6573
rect 3454 -6997 3793 -6877
rect 43568 -7728 43904 -5096
rect 8008 -7896 43904 -7728
rect 4846 -8302 5484 -8297
rect 4846 -8355 4893 -8302
rect 4956 -8355 5484 -8302
rect 4846 -8361 5484 -8355
rect 4406 -8473 5280 -8409
rect 3471 -9013 3697 -8893
rect 3656 -9317 3851 -9307
rect 3656 -9373 3696 -9317
rect 3752 -9373 3851 -9317
rect 8040 -9365 8116 -7896
rect 9713 -8301 10374 -8297
rect 9713 -8354 9772 -8301
rect 9834 -8354 10374 -8301
rect 9713 -8361 10374 -8354
rect 9230 -8473 10144 -8409
rect 3656 -9383 3851 -9373
rect 8551 -9383 8566 -9307
rect 8627 -9383 8704 -9307
rect 12886 -9365 12962 -7896
rect 14549 -8305 15056 -8297
rect 14549 -8357 14580 -8305
rect 14645 -8357 15056 -8305
rect 14549 -8361 15056 -8357
rect 14093 -8473 15025 -8409
rect 17732 -9365 17808 -7896
rect 19371 -8306 19899 -8297
rect 19371 -8358 19458 -8306
rect 19521 -8358 19899 -8306
rect 19371 -8361 19899 -8358
rect 18905 -8473 20398 -8409
rect 18241 -9321 18368 -9307
rect 18241 -9373 18256 -9321
rect 18314 -9373 18368 -9321
rect 22578 -9365 22654 -7896
rect 24212 -8303 24784 -8297
rect 24212 -8356 24269 -8303
rect 24334 -8356 24784 -8303
rect 24212 -8361 24784 -8356
rect 23789 -8473 25283 -8409
rect 27424 -9365 27500 -7896
rect 29050 -8305 29560 -8297
rect 29050 -8358 29145 -8305
rect 29206 -8358 29560 -8305
rect 29050 -8361 29560 -8358
rect 28617 -8473 30052 -8409
rect 27976 -9317 28074 -9307
rect 18241 -9383 18368 -9373
rect 27976 -9375 27993 -9317
rect 28053 -9375 28074 -9317
rect 32270 -9365 32346 -7896
rect 33926 -8305 34713 -8297
rect 33926 -8357 33989 -8305
rect 34051 -8357 34713 -8305
rect 33926 -8361 34713 -8357
rect 33465 -8473 34789 -8409
rect 32853 -9317 32953 -9307
rect 27976 -9383 28074 -9375
rect 32853 -9372 32868 -9317
rect 32932 -9372 32953 -9317
rect 37116 -9365 37192 -7896
rect 37745 -8252 37796 -8092
rect 38769 -8306 39440 -8297
rect 38769 -8358 38833 -8306
rect 38894 -8358 39440 -8306
rect 38769 -8361 39440 -8358
rect 38350 -8473 39689 -8409
rect 41962 -9365 42038 -7896
rect 32853 -9383 32953 -9372
rect 3482 -9797 3708 -9677
rect 43568 -10528 43904 -7896
rect 8008 -10696 43904 -10528
rect 3489 -10909 3772 -10789
rect 4846 -11102 5484 -11097
rect 4846 -11155 4893 -11102
rect 4956 -11155 5484 -11102
rect 4846 -11161 5484 -11155
rect 4406 -11273 5280 -11209
rect 3472 -11813 3818 -11573
rect 2863 -11970 2929 -11959
rect 3676 -12183 3688 -12107
rect 3758 -12183 3872 -12107
rect 8040 -12165 8116 -10696
rect 9713 -11101 10374 -11097
rect 9713 -11154 9772 -11101
rect 9834 -11154 10374 -11101
rect 9713 -11161 10374 -11154
rect 9230 -11273 10144 -11209
rect 8541 -12118 8702 -12107
rect 8541 -12171 8562 -12118
rect 8614 -12171 8702 -12118
rect 12886 -12165 12962 -10696
rect 14549 -11105 15056 -11097
rect 14549 -11157 14580 -11105
rect 14645 -11157 15056 -11105
rect 14549 -11161 15056 -11157
rect 14093 -11273 15025 -11209
rect 17732 -12165 17808 -10696
rect 19371 -11106 19899 -11097
rect 19371 -11158 19458 -11106
rect 19521 -11158 19899 -11106
rect 19371 -11161 19899 -11158
rect 18905 -11273 20398 -11209
rect 18239 -12121 18373 -12107
rect 8541 -12183 8702 -12171
rect 18239 -12174 18253 -12121
rect 18309 -12174 18373 -12121
rect 22578 -12165 22654 -10696
rect 24212 -11103 24784 -11097
rect 24212 -11156 24269 -11103
rect 24334 -11156 24784 -11103
rect 24212 -11161 24784 -11156
rect 23789 -11273 25283 -11209
rect 27424 -12165 27500 -10696
rect 29050 -11105 29560 -11097
rect 29050 -11158 29145 -11105
rect 29206 -11158 29560 -11105
rect 29050 -11161 29560 -11158
rect 28617 -11273 30052 -11209
rect 27983 -12117 28075 -12107
rect 18239 -12183 18373 -12174
rect 27983 -12175 27998 -12117
rect 28058 -12175 28075 -12117
rect 32270 -12165 32346 -10696
rect 33926 -11105 34788 -11097
rect 33926 -11157 33989 -11105
rect 34051 -11157 34788 -11105
rect 33926 -11161 34788 -11157
rect 33465 -11273 34789 -11209
rect 32836 -12119 32933 -12107
rect 27983 -12183 28075 -12175
rect 32836 -12171 32889 -12119
rect 37116 -12165 37192 -10696
rect 37744 -11052 37796 -10893
rect 38769 -11106 39440 -11097
rect 38769 -11158 38833 -11106
rect 38894 -11158 39440 -11106
rect 38769 -11161 39440 -11158
rect 38350 -11273 39689 -11209
rect 41962 -12165 42038 -10696
rect 32836 -12183 32933 -12171
rect 3501 -12597 3765 -12477
rect 43568 -13328 43904 -10696
rect 8008 -13496 43904 -13328
rect 4846 -13902 5484 -13897
rect 4846 -13955 4893 -13902
rect 4956 -13955 5484 -13902
rect 4846 -13961 5484 -13955
rect 4406 -14073 5280 -14009
rect 3478 -14613 3710 -14493
rect 3668 -14983 3681 -14907
rect 3746 -14983 3864 -14907
rect 8040 -14965 8116 -13496
rect 9713 -13901 10374 -13897
rect 9713 -13954 9772 -13901
rect 9834 -13954 10374 -13901
rect 9713 -13961 10374 -13954
rect 9230 -14073 10144 -14009
rect 8561 -14919 8697 -14907
rect 8561 -14971 8581 -14919
rect 8633 -14971 8697 -14919
rect 12886 -14965 12962 -13496
rect 14549 -13905 15056 -13897
rect 14549 -13957 14580 -13905
rect 14645 -13957 15056 -13905
rect 14549 -13961 15056 -13957
rect 14093 -14073 15025 -14009
rect 17732 -14965 17808 -13496
rect 19371 -13906 19899 -13897
rect 19371 -13958 19458 -13906
rect 19521 -13958 19899 -13906
rect 19371 -13961 19899 -13958
rect 18905 -14073 20398 -14009
rect 18243 -14921 18383 -14907
rect 8561 -14983 8697 -14971
rect 18243 -14974 18256 -14921
rect 18312 -14974 18383 -14921
rect 22578 -14965 22654 -13496
rect 24212 -13903 24784 -13897
rect 24212 -13956 24269 -13903
rect 24334 -13956 24784 -13903
rect 24212 -13961 24784 -13956
rect 23789 -14073 25283 -14009
rect 27424 -14965 27500 -13496
rect 29050 -13905 29560 -13897
rect 29050 -13958 29145 -13905
rect 29206 -13958 29560 -13905
rect 29050 -13961 29560 -13958
rect 28617 -14073 30052 -14009
rect 27977 -14916 28064 -14907
rect 18243 -14983 18383 -14974
rect 27977 -14972 27997 -14916
rect 28062 -14972 28064 -14916
rect 32270 -14965 32346 -13496
rect 33926 -13905 34722 -13897
rect 33926 -13957 33989 -13905
rect 34051 -13957 34722 -13905
rect 33926 -13961 34722 -13957
rect 33465 -14073 34789 -14009
rect 32847 -14918 32968 -14907
rect 27977 -14983 28064 -14972
rect 32847 -14973 32868 -14918
rect 32936 -14973 32968 -14918
rect 37116 -14965 37192 -13496
rect 37751 -13709 37796 -13704
rect 37750 -13852 37796 -13709
rect 38769 -13906 39440 -13897
rect 38769 -13958 38833 -13906
rect 38894 -13958 39440 -13906
rect 38769 -13961 39440 -13958
rect 38350 -14073 39689 -14009
rect 41962 -14965 42038 -13496
rect 32847 -14983 32968 -14973
rect 3480 -15397 3712 -15277
rect 43568 -16128 43904 -13496
rect 8008 -16296 43904 -16128
rect 3473 -16509 3739 -16389
rect 4846 -16702 5484 -16697
rect 4846 -16755 4893 -16702
rect 4956 -16755 5484 -16702
rect 4846 -16761 5484 -16755
rect 4406 -16873 5280 -16809
rect 3455 -17413 3722 -17173
rect 3674 -17783 3692 -17707
rect 3760 -17783 3881 -17707
rect 8040 -17765 8116 -16296
rect 9713 -16701 10374 -16697
rect 9713 -16754 9772 -16701
rect 9834 -16754 10374 -16701
rect 9713 -16761 10374 -16754
rect 9230 -16873 10144 -16809
rect 8551 -17720 8709 -17707
rect 8551 -17772 8572 -17720
rect 8626 -17772 8709 -17720
rect 12886 -17765 12962 -16296
rect 14549 -16705 15056 -16697
rect 14549 -16757 14580 -16705
rect 14645 -16757 15056 -16705
rect 14549 -16761 15056 -16757
rect 14093 -16873 15025 -16809
rect 17732 -17765 17808 -16296
rect 19371 -16706 19899 -16697
rect 19371 -16758 19458 -16706
rect 19521 -16758 19899 -16706
rect 19371 -16761 19899 -16758
rect 18905 -16873 20398 -16809
rect 18239 -17717 18381 -17707
rect 8551 -17783 8709 -17772
rect 18239 -17773 18253 -17717
rect 18315 -17773 18381 -17717
rect 22578 -17765 22654 -16296
rect 24212 -16703 24784 -16697
rect 24212 -16756 24269 -16703
rect 24334 -16756 24784 -16703
rect 24212 -16761 24784 -16756
rect 23789 -16873 25283 -16809
rect 18239 -17783 18381 -17773
rect 27424 -17765 27500 -16296
rect 29050 -16705 29560 -16697
rect 29050 -16758 29145 -16705
rect 29206 -16758 29560 -16705
rect 29050 -16761 29560 -16758
rect 28617 -16873 30052 -16809
rect 27987 -17716 28062 -17707
rect 27987 -17769 27999 -17716
rect 28060 -17769 28062 -17716
rect 32270 -17765 32346 -16296
rect 33926 -16705 34695 -16697
rect 33926 -16757 33989 -16705
rect 34051 -16757 34695 -16705
rect 33926 -16761 34695 -16757
rect 33465 -16873 34789 -16809
rect 32842 -17715 32947 -17707
rect 27987 -17783 28062 -17769
rect 32842 -17775 32868 -17715
rect 32935 -17775 32947 -17715
rect 37116 -17765 37192 -16296
rect 38769 -16706 39440 -16697
rect 38769 -16758 38833 -16706
rect 38894 -16758 39440 -16706
rect 38769 -16761 39440 -16758
rect 38350 -16873 39689 -16809
rect 41962 -17765 42038 -16296
rect 32842 -17783 32947 -17775
rect 3477 -18197 3695 -18077
rect 38732 -18928 38984 -18927
rect 43568 -18928 43904 -16296
rect 8008 -19096 43904 -18928
rect 3824 -19452 3874 -19286
rect 4846 -19502 5484 -19497
rect 4846 -19555 4893 -19502
rect 4956 -19555 5484 -19502
rect 4846 -19561 5484 -19555
rect 4406 -19673 5280 -19609
rect 3679 -20583 3696 -20507
rect 3752 -20583 3853 -20507
rect 8040 -20565 8116 -19096
rect 8670 -19452 8720 -19286
rect 9713 -19501 10374 -19497
rect 9713 -19554 9772 -19501
rect 9834 -19554 10374 -19501
rect 9713 -19561 10374 -19554
rect 9230 -19673 10144 -19609
rect 8557 -20518 8706 -20507
rect 8557 -20570 8568 -20518
rect 8620 -20570 8706 -20518
rect 12886 -20565 12962 -19096
rect 13516 -19452 13566 -19286
rect 14549 -19505 15056 -19497
rect 14549 -19557 14580 -19505
rect 14645 -19557 15056 -19505
rect 14549 -19561 15056 -19557
rect 14093 -19673 15025 -19609
rect 17732 -20565 17808 -19096
rect 18362 -19452 18412 -19286
rect 19371 -19506 19899 -19497
rect 19371 -19558 19458 -19506
rect 19521 -19558 19899 -19506
rect 19371 -19561 19899 -19558
rect 18905 -19673 20398 -19609
rect 18239 -20521 18374 -20507
rect 8557 -20583 8706 -20570
rect 18239 -20577 18254 -20521
rect 18312 -20577 18374 -20521
rect 22578 -20565 22654 -19096
rect 23208 -19452 23258 -19286
rect 24212 -19503 24784 -19497
rect 24212 -19556 24269 -19503
rect 24334 -19556 24784 -19503
rect 24212 -19561 24784 -19556
rect 23789 -19673 25283 -19609
rect 27424 -20565 27500 -19096
rect 28054 -19452 28104 -19286
rect 29050 -19505 29560 -19497
rect 29050 -19558 29145 -19505
rect 29206 -19558 29560 -19505
rect 29050 -19561 29560 -19558
rect 28617 -19673 30052 -19609
rect 27988 -20517 28074 -20507
rect 27988 -20574 27998 -20517
rect 28059 -20574 28074 -20517
rect 32270 -20565 32346 -19096
rect 32900 -19452 32950 -19286
rect 33926 -19505 35419 -19497
rect 33926 -19557 33989 -19505
rect 34051 -19557 35419 -19505
rect 33926 -19561 35419 -19557
rect 33465 -19673 34789 -19609
rect 32844 -20517 32953 -20507
rect 18239 -20583 18374 -20577
rect 27988 -20583 28074 -20574
rect 32844 -20574 32869 -20517
rect 32932 -20574 32953 -20517
rect 37116 -20565 37192 -19096
rect 43568 -19219 43904 -19096
rect 32844 -20583 32953 -20574
<< via1 >>
rect 3696 2436 3752 2492
rect 8568 2436 8624 2492
rect 13496 2438 13552 2494
rect 18256 2435 18312 2491
rect 23184 2436 23240 2492
rect 28000 2441 28056 2497
rect 32872 2408 32928 2464
rect 3107 1757 3167 1818
rect 13719 1206 13776 1273
rect 18565 1188 18626 1254
rect 23407 1229 23464 1298
rect 28280 1224 28337 1287
rect 33095 1202 33156 1262
rect 2765 836 2823 890
rect 6722 822 6785 883
rect 4032 485 4088 537
rect 3802 -93 3874 -37
rect 4035 -67 4089 -15
rect 3107 -314 3167 -197
rect 2769 -776 2822 -683
rect 3112 -977 3165 -924
rect 3700 -983 3768 -907
rect 7569 -952 7623 -899
rect 8648 -93 8720 -36
rect 8882 -66 8934 -14
rect 8574 -983 8632 -907
rect 12415 -952 12469 -899
rect 13494 -93 13566 -38
rect 13727 -67 13782 -15
rect 13505 -974 13567 -916
rect 17261 -952 17315 -899
rect 18340 -90 18412 -34
rect 18573 -68 18628 -15
rect 18259 -970 18311 -918
rect 22107 -952 22161 -899
rect 23186 -88 23258 -33
rect 23420 -67 23474 -14
rect 23199 -968 23256 -916
rect 26953 -952 27007 -899
rect 28032 -89 28104 -34
rect 28264 -67 28322 -15
rect 28001 -971 28056 -918
rect 31799 -952 31853 -899
rect 32878 -91 32950 -35
rect 33111 -68 33166 -15
rect 32869 -972 32932 -915
rect 36645 -952 36699 -899
rect 37959 -66 38011 -14
rect 41491 -952 41545 -899
rect 7602 -1104 7656 -1051
rect 8019 -1103 8073 -1050
rect 12448 -1104 12502 -1051
rect 12865 -1103 12919 -1050
rect 17294 -1104 17348 -1051
rect 17711 -1103 17765 -1050
rect 22140 -1104 22194 -1051
rect 22557 -1103 22611 -1050
rect 26986 -1104 27040 -1051
rect 27403 -1103 27457 -1050
rect 31832 -1104 31886 -1051
rect 32249 -1103 32303 -1050
rect 36678 -1104 36732 -1051
rect 37095 -1103 37149 -1050
rect 41524 -1104 41578 -1051
rect 41941 -1103 41995 -1050
rect 4893 -2755 4956 -2702
rect 3802 -2891 3874 -2835
rect 4037 -2867 4090 -2814
rect 3095 -3778 3148 -3721
rect 3687 -3783 3755 -3707
rect 7569 -3752 7623 -3699
rect 9772 -2754 9834 -2701
rect 8648 -2893 8720 -2837
rect 8882 -2867 8936 -2815
rect 8568 -3783 8628 -3707
rect 12415 -3752 12469 -3699
rect 14580 -2757 14645 -2705
rect 13494 -2892 13566 -2835
rect 13727 -2867 13782 -2814
rect 13510 -3772 13566 -3717
rect 17261 -3752 17315 -3699
rect 19458 -2758 19521 -2706
rect 18340 -2891 18412 -2835
rect 18573 -2867 18627 -2815
rect 18261 -3773 18319 -3719
rect 22107 -3752 22161 -3699
rect 24269 -2756 24334 -2703
rect 23186 -2890 23258 -2834
rect 23418 -2868 23472 -2815
rect 23194 -3774 23253 -3718
rect 26953 -3752 27007 -3699
rect 29145 -2758 29206 -2705
rect 28032 -2890 28104 -2834
rect 28267 -2866 28320 -2812
rect 27993 -3770 28049 -3718
rect 31799 -3752 31853 -3699
rect 33989 -2757 34051 -2705
rect 32878 -2889 32950 -2832
rect 33112 -2867 33164 -2815
rect 32869 -3774 32932 -3714
rect 36645 -3752 36699 -3699
rect 38833 -2758 38894 -2706
rect 37724 -2892 37796 -2834
rect 41491 -3752 41545 -3699
rect 7602 -3904 7656 -3851
rect 8019 -3903 8073 -3850
rect 12448 -3904 12502 -3851
rect 12865 -3903 12919 -3850
rect 17294 -3904 17348 -3851
rect 17711 -3903 17765 -3850
rect 22140 -3904 22194 -3851
rect 22557 -3903 22611 -3850
rect 26986 -3904 27040 -3851
rect 27403 -3903 27457 -3850
rect 31832 -3904 31886 -3851
rect 32249 -3903 32303 -3850
rect 36678 -3904 36732 -3851
rect 37095 -3903 37149 -3850
rect 41524 -3904 41578 -3851
rect 41941 -3903 41995 -3850
rect 4893 -5555 4956 -5502
rect 3802 -5693 3874 -5637
rect 4037 -5666 4089 -5614
rect 3076 -5907 3146 -5826
rect 2750 -6351 2803 -6277
rect 3091 -6566 3143 -6514
rect 3691 -6583 3750 -6507
rect 7569 -6552 7623 -6499
rect 9772 -5554 9834 -5501
rect 8648 -5690 8720 -5632
rect 8882 -5667 8935 -5615
rect 8565 -6583 8624 -6507
rect 12415 -6552 12469 -6499
rect 14580 -5557 14645 -5505
rect 13494 -5692 13566 -5635
rect 13728 -5667 13780 -5615
rect 13508 -6571 13566 -6515
rect 17261 -6552 17315 -6499
rect 19458 -5558 19521 -5506
rect 18340 -5691 18412 -5634
rect 18574 -5667 18629 -5612
rect 18257 -6573 18315 -6520
rect 22107 -6552 22161 -6499
rect 24269 -5556 24334 -5503
rect 23186 -5691 23258 -5634
rect 23420 -5667 23473 -5614
rect 23194 -6572 23250 -6517
rect 26953 -6552 27007 -6499
rect 29145 -5558 29206 -5505
rect 28032 -5691 28104 -5634
rect 28267 -5666 28319 -5614
rect 27989 -6574 28042 -6519
rect 31799 -6552 31853 -6499
rect 33989 -5557 34051 -5505
rect 32878 -5691 32950 -5634
rect 33111 -5667 33165 -5614
rect 32870 -6573 32933 -6518
rect 36645 -6552 36699 -6499
rect 38833 -5558 38894 -5506
rect 37959 -5666 38011 -5614
rect 41491 -6552 41545 -6499
rect 7602 -6704 7656 -6651
rect 8019 -6703 8073 -6650
rect 12448 -6704 12502 -6651
rect 12865 -6703 12919 -6650
rect 17294 -6704 17348 -6651
rect 17711 -6703 17765 -6650
rect 22140 -6704 22194 -6651
rect 22557 -6703 22611 -6650
rect 26986 -6704 27040 -6651
rect 27403 -6703 27457 -6650
rect 31832 -6704 31886 -6651
rect 32249 -6703 32303 -6650
rect 36678 -6704 36732 -6651
rect 37095 -6703 37149 -6650
rect 41524 -6704 41578 -6651
rect 41941 -6703 41995 -6650
rect 4893 -8355 4956 -8302
rect 3802 -8493 3874 -8434
rect 4036 -8467 4089 -8415
rect 3696 -9373 3752 -9317
rect 7569 -9352 7623 -9299
rect 9772 -8354 9834 -8301
rect 8648 -8492 8720 -8435
rect 8882 -8469 8938 -8414
rect 8566 -9383 8627 -9307
rect 12415 -9352 12469 -9299
rect 14580 -8357 14645 -8305
rect 13494 -8491 13566 -8433
rect 13728 -8467 13780 -8415
rect 13510 -9371 13567 -9316
rect 17261 -9352 17315 -9299
rect 19458 -8358 19521 -8306
rect 18340 -8491 18412 -8433
rect 18571 -8470 18629 -8412
rect 18256 -9373 18314 -9321
rect 22107 -9352 22161 -9299
rect 24269 -8356 24334 -8303
rect 23186 -8491 23258 -8434
rect 23420 -8468 23475 -8413
rect 23196 -9371 23250 -9316
rect 26953 -9352 27007 -9299
rect 29145 -8358 29206 -8305
rect 28032 -8492 28104 -8433
rect 28264 -8467 28321 -8413
rect 27993 -9375 28053 -9317
rect 31799 -9352 31853 -9299
rect 33989 -8357 34051 -8305
rect 32878 -8490 32950 -8434
rect 33110 -8469 33165 -8414
rect 32868 -9372 32932 -9317
rect 36645 -9352 36699 -9299
rect 38833 -8358 38894 -8306
rect 37958 -8467 38010 -8415
rect 41491 -9352 41545 -9299
rect 3298 -9464 3362 -9400
rect 7602 -9504 7656 -9451
rect 8019 -9503 8073 -9450
rect 12448 -9504 12502 -9451
rect 12865 -9503 12919 -9450
rect 17294 -9504 17348 -9451
rect 17711 -9503 17765 -9450
rect 22140 -9504 22194 -9451
rect 22557 -9503 22611 -9450
rect 26986 -9504 27040 -9451
rect 27403 -9503 27457 -9450
rect 31832 -9504 31886 -9451
rect 32249 -9503 32303 -9450
rect 36678 -9504 36732 -9451
rect 37095 -9503 37149 -9450
rect 41524 -9504 41578 -9451
rect 41941 -9503 41995 -9450
rect 4893 -11155 4956 -11102
rect 3802 -11291 3874 -11232
rect 4037 -11266 4089 -11214
rect 3096 -11514 3157 -11421
rect 2865 -11959 2926 -11876
rect 3202 -12225 3262 -12159
rect 3688 -12183 3758 -12107
rect 7569 -12152 7623 -12099
rect 9772 -11154 9834 -11101
rect 8648 -11291 8720 -11235
rect 8874 -11272 8938 -11212
rect 8562 -12171 8614 -12118
rect 12415 -12152 12469 -12099
rect 14580 -11157 14645 -11105
rect 13494 -11293 13566 -11233
rect 13728 -11266 13780 -11214
rect 13506 -12171 13560 -12119
rect 17261 -12152 17315 -12099
rect 19458 -11158 19521 -11106
rect 18340 -11291 18412 -11231
rect 18573 -11268 18626 -11213
rect 18253 -12174 18309 -12121
rect 22107 -12152 22161 -12099
rect 24269 -11156 24334 -11103
rect 23186 -11293 23258 -11235
rect 23420 -11267 23477 -11213
rect 23192 -12173 23252 -12116
rect 26953 -12152 27007 -12099
rect 29145 -11158 29206 -11105
rect 28032 -11291 28104 -11234
rect 28266 -11266 28318 -11214
rect 27998 -12175 28058 -12117
rect 31799 -12152 31853 -12099
rect 33989 -11157 34051 -11105
rect 32878 -11291 32950 -11234
rect 33111 -11268 33164 -11216
rect 32889 -12171 32941 -12119
rect 36645 -12152 36699 -12099
rect 38833 -11158 38894 -11106
rect 37956 -11269 38014 -11213
rect 41491 -12152 41545 -12099
rect 7602 -12304 7656 -12251
rect 8019 -12303 8073 -12250
rect 12448 -12304 12502 -12251
rect 12865 -12303 12919 -12250
rect 17294 -12304 17348 -12251
rect 17711 -12303 17765 -12250
rect 22140 -12304 22194 -12251
rect 22557 -12303 22611 -12250
rect 26986 -12304 27040 -12251
rect 27403 -12303 27457 -12250
rect 31832 -12304 31886 -12251
rect 32249 -12303 32303 -12250
rect 36678 -12304 36732 -12251
rect 37095 -12303 37149 -12250
rect 41524 -12304 41578 -12251
rect 41941 -12303 41995 -12250
rect 4893 -13955 4956 -13902
rect 3802 -14091 3874 -14035
rect 4037 -14067 4089 -14015
rect 3185 -14976 3254 -14908
rect 3681 -14983 3746 -14907
rect 7569 -14952 7623 -14899
rect 9772 -13954 9834 -13901
rect 8648 -14091 8720 -14035
rect 8882 -14067 8937 -14013
rect 8581 -14971 8633 -14919
rect 12415 -14952 12469 -14899
rect 14580 -13957 14645 -13905
rect 13494 -14092 13566 -14035
rect 13727 -14067 13782 -14014
rect 13512 -14971 13567 -14918
rect 17261 -14952 17315 -14899
rect 19458 -13958 19521 -13906
rect 18340 -14090 18412 -14033
rect 18572 -14068 18630 -14013
rect 18256 -14974 18312 -14921
rect 22107 -14952 22161 -14899
rect 24269 -13956 24334 -13903
rect 23186 -14092 23258 -14036
rect 23419 -14068 23474 -14015
rect 23196 -14971 23251 -14913
rect 26953 -14952 27007 -14899
rect 29145 -13958 29206 -13905
rect 28032 -14093 28104 -14037
rect 28264 -14067 28320 -14013
rect 27997 -14972 28062 -14916
rect 31799 -14952 31853 -14899
rect 33989 -13957 34051 -13905
rect 32878 -14093 32950 -14037
rect 33112 -14067 33164 -14014
rect 32868 -14973 32936 -14918
rect 36645 -14952 36699 -14899
rect 38833 -13958 38894 -13906
rect 37953 -14068 38013 -14012
rect 41491 -14952 41545 -14899
rect 7602 -15104 7656 -15051
rect 8019 -15103 8073 -15050
rect 12448 -15104 12502 -15051
rect 12865 -15103 12919 -15050
rect 17294 -15104 17348 -15051
rect 17711 -15103 17765 -15050
rect 22140 -15104 22194 -15051
rect 22557 -15103 22611 -15050
rect 26986 -15104 27040 -15051
rect 27403 -15103 27457 -15050
rect 31832 -15104 31886 -15051
rect 32249 -15103 32303 -15050
rect 36678 -15104 36732 -15051
rect 37095 -15103 37149 -15050
rect 41524 -15104 41578 -15051
rect 41941 -15103 41995 -15050
rect 4893 -16755 4956 -16702
rect 3181 -16883 3251 -16806
rect 3802 -16891 3874 -16835
rect 4036 -16867 4088 -16815
rect 2850 -17778 2911 -17716
rect 3692 -17783 3760 -17707
rect 7569 -17752 7623 -17699
rect 9772 -16754 9834 -16701
rect 8648 -16892 8720 -16836
rect 8882 -16867 8934 -16815
rect 8572 -17772 8626 -17720
rect 12415 -17752 12469 -17699
rect 14580 -16757 14645 -16705
rect 13494 -16891 13566 -16835
rect 13728 -16867 13783 -16814
rect 13507 -17769 13559 -17717
rect 17261 -17752 17315 -17699
rect 19458 -16758 19521 -16706
rect 18340 -16892 18412 -16836
rect 18573 -16868 18627 -16814
rect 18253 -17773 18315 -17717
rect 22107 -17752 22161 -17699
rect 24269 -16756 24334 -16703
rect 23186 -16893 23258 -16837
rect 23419 -16867 23475 -16814
rect 23197 -17775 23250 -17714
rect 26953 -17752 27007 -17699
rect 29145 -16758 29206 -16705
rect 28032 -16893 28104 -16837
rect 28267 -16866 28320 -16814
rect 27999 -17769 28060 -17716
rect 31799 -17752 31853 -17699
rect 33989 -16757 34051 -16705
rect 32878 -16893 32950 -16835
rect 33112 -16867 33165 -16815
rect 32868 -17775 32935 -17715
rect 36645 -17752 36699 -17699
rect 38833 -16758 38894 -16706
rect 37953 -16870 38015 -16808
rect 41491 -17752 41545 -17699
rect 7602 -17904 7656 -17851
rect 8019 -17903 8073 -17850
rect 12448 -17904 12502 -17851
rect 12865 -17903 12919 -17850
rect 17294 -17904 17348 -17851
rect 17711 -17903 17765 -17850
rect 22140 -17904 22194 -17851
rect 22557 -17903 22611 -17850
rect 26986 -17904 27040 -17851
rect 27403 -17903 27457 -17850
rect 31832 -17904 31886 -17851
rect 32249 -17903 32303 -17850
rect 36678 -17904 36732 -17851
rect 37095 -17903 37149 -17850
rect 41524 -17904 41578 -17851
rect 41941 -17903 41995 -17850
rect 4893 -19555 4956 -19502
rect 4036 -19668 4089 -19615
rect 3696 -20583 3752 -20507
rect 7569 -20552 7623 -20499
rect 9772 -19554 9834 -19501
rect 8882 -19666 8936 -19614
rect 8568 -20570 8620 -20518
rect 12415 -20552 12469 -20499
rect 14580 -19557 14645 -19505
rect 13729 -19666 13781 -19614
rect 13515 -20570 13568 -20518
rect 17261 -20552 17315 -20499
rect 19458 -19558 19521 -19506
rect 18573 -19669 18630 -19613
rect 18254 -20577 18312 -20521
rect 22107 -20552 22161 -20499
rect 24269 -19556 24334 -19503
rect 23419 -19667 23474 -19615
rect 23198 -20574 23250 -20517
rect 26953 -20552 27007 -20499
rect 29145 -19558 29206 -19505
rect 28263 -19667 28318 -19614
rect 27998 -20574 28059 -20517
rect 31799 -20552 31853 -20499
rect 33989 -19557 34051 -19505
rect 33111 -19668 33166 -19614
rect 32869 -20574 32932 -20517
rect 36645 -20552 36699 -20499
rect 7602 -20704 7656 -20651
rect 8019 -20703 8073 -20650
rect 12448 -20704 12502 -20651
rect 12865 -20703 12919 -20650
rect 17294 -20704 17348 -20651
rect 17711 -20703 17765 -20650
rect 22140 -20704 22194 -20651
rect 22557 -20703 22611 -20650
rect 26986 -20704 27040 -20651
rect 27403 -20703 27457 -20650
rect 31832 -20704 31886 -20651
rect 32249 -20703 32303 -20650
rect 36678 -20704 36732 -20651
rect 37095 -20703 37149 -20650
<< metal2 >>
rect 3686 2492 3762 2502
rect 3686 2436 3696 2492
rect 3752 2436 3762 2492
rect 3686 2426 3762 2436
rect 8558 2492 8634 2502
rect 8558 2436 8568 2492
rect 8624 2436 8634 2492
rect 8558 2426 8634 2436
rect 13486 2494 13562 2504
rect 13486 2438 13496 2494
rect 13552 2438 13562 2494
rect 13486 2428 13562 2438
rect 18246 2491 18322 2501
rect 18246 2435 18256 2491
rect 18312 2435 18322 2491
rect 18246 2425 18322 2435
rect 23174 2492 23250 2502
rect 23174 2436 23184 2492
rect 23240 2436 23250 2492
rect 23174 2426 23250 2436
rect 27987 2497 28069 2509
rect 27987 2441 28000 2497
rect 28056 2441 28069 2497
rect 27987 2429 28069 2441
rect 32858 2464 32939 2476
rect 32858 2408 32872 2464
rect 32928 2408 32939 2464
rect 32858 2394 32939 2408
rect 3089 1818 3185 1835
rect 3089 1757 3107 1818
rect 3167 1757 3185 1818
rect 3089 1736 3185 1757
rect 2749 890 2835 897
rect 2749 836 2765 890
rect 2823 889 2835 890
rect 3101 889 3169 1736
rect 23370 1301 23497 1314
rect 13688 1278 13804 1299
rect 13688 1203 13716 1278
rect 13780 1203 13804 1278
rect 13688 1181 13804 1203
rect 18536 1257 18648 1264
rect 18536 1185 18562 1257
rect 18631 1185 18648 1257
rect 23370 1223 23403 1301
rect 23468 1223 23497 1301
rect 23370 1196 23497 1223
rect 28247 1291 28370 1304
rect 28247 1218 28271 1291
rect 28344 1218 28370 1291
rect 28247 1192 28370 1218
rect 33065 1262 33188 1274
rect 33065 1202 33095 1262
rect 33156 1202 33188 1262
rect 18536 1166 18648 1185
rect 33065 1176 33188 1202
rect 43064 896 43400 1400
rect 2823 836 3170 889
rect 2749 821 3170 836
rect 6693 888 6807 894
rect 6693 819 6718 888
rect 6790 819 6807 888
rect 6693 804 6807 819
rect 7504 728 43400 896
rect 3998 537 4115 539
rect 3998 480 4029 537
rect 4093 480 4115 537
rect 3998 448 4115 480
rect 4010 -13 4115 -1
rect 3782 -37 3919 -28
rect 3782 -93 3802 -37
rect 3874 -93 3919 -37
rect 4010 -69 4033 -13
rect 4092 -69 4115 -13
rect 4010 -78 4115 -69
rect 3782 -105 3919 -93
rect 3099 -197 3170 -163
rect 3099 -255 3107 -197
rect 2759 -314 3107 -255
rect 3167 -314 3170 -197
rect 2759 -327 3170 -314
rect 2759 -683 2831 -327
rect 2759 -776 2769 -683
rect 2822 -776 2831 -683
rect 2759 -800 2831 -776
rect 3098 -922 3174 -897
rect 3098 -980 3110 -922
rect 3168 -980 3174 -922
rect 3098 -1001 3174 -980
rect 3672 -907 3794 -884
rect 3672 -983 3696 -907
rect 3774 -983 3794 -907
rect 7558 -899 7634 728
rect 8859 -12 8951 -8
rect 8624 -36 8758 -27
rect 8624 -93 8648 -36
rect 8720 -93 8758 -36
rect 8859 -68 8880 -12
rect 8938 -68 8951 -12
rect 8859 -74 8951 -68
rect 8624 -103 8758 -93
rect 7558 -952 7569 -899
rect 7623 -952 7634 -899
rect 7558 -965 7634 -952
rect 8545 -907 8658 -893
rect 3672 -1002 3794 -983
rect 8545 -983 8574 -907
rect 8632 -983 8658 -907
rect 12404 -899 12480 728
rect 13701 -13 13810 -1
rect 13466 -37 13600 -29
rect 13466 -93 13494 -37
rect 13566 -93 13600 -37
rect 13701 -69 13725 -13
rect 13784 -69 13810 -13
rect 13701 -78 13810 -69
rect 13466 -105 13600 -93
rect 12404 -952 12415 -899
rect 12469 -952 12480 -899
rect 12404 -965 12480 -952
rect 13469 -916 13581 -896
rect 8545 -1000 8658 -983
rect 13469 -974 13505 -916
rect 13567 -974 13581 -916
rect 17250 -899 17326 728
rect 18553 -12 18646 2
rect 18312 -34 18442 -29
rect 18312 -90 18340 -34
rect 18412 -90 18442 -34
rect 18553 -70 18570 -12
rect 18632 -70 18646 -12
rect 18553 -84 18646 -70
rect 18312 -105 18442 -90
rect 17250 -952 17261 -899
rect 17315 -952 17326 -899
rect 17250 -965 17326 -952
rect 18223 -915 18325 -896
rect 13469 -998 13581 -974
rect 18223 -972 18256 -915
rect 18315 -972 18325 -915
rect 22096 -899 22172 728
rect 23405 -12 23487 -1
rect 23154 -32 23295 -29
rect 23154 -88 23186 -32
rect 23258 -88 23295 -32
rect 23405 -69 23418 -12
rect 23476 -69 23487 -12
rect 23405 -80 23487 -69
rect 23154 -105 23295 -88
rect 22096 -952 22107 -899
rect 22161 -952 22172 -899
rect 22096 -965 22172 -952
rect 23156 -913 23270 -895
rect 18223 -996 18325 -972
rect 23156 -971 23194 -913
rect 23260 -971 23270 -913
rect 26942 -899 27018 728
rect 28249 -13 28338 1
rect 28000 -33 28138 -29
rect 28000 -89 28032 -33
rect 28104 -89 28138 -33
rect 28249 -69 28262 -13
rect 28325 -69 28338 -13
rect 28249 -83 28338 -69
rect 28000 -105 28138 -89
rect 26942 -952 26953 -899
rect 27007 -952 27018 -899
rect 26942 -965 27018 -952
rect 27975 -915 28081 -898
rect 23156 -999 23270 -971
rect 27975 -975 27999 -915
rect 28058 -975 28081 -915
rect 31788 -899 31864 728
rect 33097 -13 33182 -3
rect 32853 -35 32979 -29
rect 32853 -91 32878 -35
rect 32950 -91 32979 -35
rect 33097 -70 33109 -13
rect 33168 -70 33182 -13
rect 33097 -79 33182 -70
rect 32853 -105 32979 -91
rect 31788 -952 31799 -899
rect 31853 -952 31864 -899
rect 31788 -965 31864 -952
rect 32850 -915 32947 -897
rect 27975 -1001 28081 -975
rect 32850 -972 32869 -915
rect 32932 -972 32947 -915
rect 36634 -899 36710 728
rect 37941 -13 38025 -4
rect 37941 -69 37955 -13
rect 38012 -69 38025 -13
rect 37941 -79 38025 -69
rect 36634 -952 36645 -899
rect 36699 -952 36710 -899
rect 36634 -965 36710 -952
rect 41480 -899 41556 728
rect 41480 -952 41491 -899
rect 41545 -952 41556 -899
rect 41480 -965 41556 -952
rect 32850 -990 32947 -972
rect 7591 -1050 8083 -1039
rect 7591 -1051 8019 -1050
rect 7591 -1104 7602 -1051
rect 7656 -1103 8019 -1051
rect 8073 -1103 8083 -1050
rect 7656 -1104 8083 -1103
rect 7591 -1115 8083 -1104
rect 12437 -1050 12929 -1039
rect 12437 -1051 12865 -1050
rect 12437 -1104 12448 -1051
rect 12502 -1103 12865 -1051
rect 12919 -1103 12929 -1050
rect 12502 -1104 12929 -1103
rect 12437 -1115 12929 -1104
rect 17283 -1050 17775 -1039
rect 17283 -1051 17711 -1050
rect 17283 -1104 17294 -1051
rect 17348 -1103 17711 -1051
rect 17765 -1103 17775 -1050
rect 17348 -1104 17775 -1103
rect 17283 -1115 17775 -1104
rect 22129 -1050 22621 -1039
rect 22129 -1051 22557 -1050
rect 22129 -1104 22140 -1051
rect 22194 -1103 22557 -1051
rect 22611 -1103 22621 -1050
rect 22194 -1104 22621 -1103
rect 22129 -1115 22621 -1104
rect 26975 -1050 27467 -1039
rect 26975 -1051 27403 -1050
rect 26975 -1104 26986 -1051
rect 27040 -1103 27403 -1051
rect 27457 -1103 27467 -1050
rect 27040 -1104 27467 -1103
rect 26975 -1115 27467 -1104
rect 31821 -1050 32313 -1039
rect 31821 -1051 32249 -1050
rect 31821 -1104 31832 -1051
rect 31886 -1103 32249 -1051
rect 32303 -1103 32313 -1050
rect 31886 -1104 32313 -1103
rect 31821 -1115 32313 -1104
rect 36667 -1050 37159 -1039
rect 36667 -1051 37095 -1050
rect 36667 -1104 36678 -1051
rect 36732 -1103 37095 -1051
rect 37149 -1103 37159 -1050
rect 36732 -1104 37159 -1103
rect 36667 -1115 37159 -1104
rect 41513 -1050 42005 -1039
rect 41513 -1051 41941 -1050
rect 41513 -1104 41524 -1051
rect 41578 -1103 41941 -1051
rect 41995 -1103 42005 -1050
rect 41578 -1104 42005 -1103
rect 41513 -1115 42005 -1104
rect 7798 -1456 7874 -1115
rect 12644 -1456 12720 -1115
rect 17490 -1456 17566 -1115
rect 22336 -1456 22412 -1115
rect 27182 -1456 27258 -1115
rect 32028 -1456 32104 -1115
rect 36874 -1456 36950 -1115
rect 41720 -1456 41796 -1115
rect 7392 -1624 42616 -1456
rect 42784 -1624 42852 -1456
rect 43064 -1904 43400 728
rect 7504 -2072 43400 -1904
rect 4872 -2699 4984 -2697
rect 4872 -2755 4893 -2699
rect 4956 -2755 4984 -2699
rect 4872 -2761 4984 -2755
rect 4009 -2812 4115 -2806
rect 3768 -2835 3902 -2828
rect 3768 -2891 3802 -2835
rect 3874 -2891 3902 -2835
rect 4009 -2868 4035 -2812
rect 4092 -2868 4115 -2812
rect 4009 -2875 4115 -2868
rect 3768 -2905 3902 -2891
rect 3082 -3720 3158 -3702
rect 3082 -3780 3092 -3720
rect 3151 -3780 3158 -3720
rect 3082 -3798 3158 -3780
rect 3655 -3707 3779 -3692
rect 3655 -3783 3687 -3707
rect 3755 -3783 3779 -3707
rect 7558 -3699 7634 -2072
rect 9744 -2698 9856 -2697
rect 9744 -2754 9772 -2698
rect 9834 -2754 9856 -2698
rect 9744 -2761 9856 -2754
rect 8860 -2812 8959 -2807
rect 8624 -2837 8748 -2828
rect 8624 -2893 8648 -2837
rect 8720 -2893 8748 -2837
rect 8860 -2870 8879 -2812
rect 8938 -2870 8959 -2812
rect 8860 -2876 8959 -2870
rect 8624 -2905 8748 -2893
rect 7558 -3752 7569 -3699
rect 7623 -3752 7634 -3699
rect 7558 -3765 7634 -3752
rect 8539 -3707 8643 -3693
rect 3655 -3800 3779 -3783
rect 8539 -3783 8568 -3707
rect 8628 -3783 8643 -3707
rect 12404 -3699 12480 -2072
rect 14560 -2701 14672 -2697
rect 14560 -2757 14580 -2701
rect 14645 -2757 14672 -2701
rect 14560 -2761 14672 -2757
rect 13704 -2812 13805 -2804
rect 13469 -2835 13590 -2828
rect 13469 -2892 13494 -2835
rect 13566 -2892 13590 -2835
rect 13704 -2869 13725 -2812
rect 13784 -2869 13805 -2812
rect 13704 -2882 13805 -2869
rect 13469 -2905 13590 -2892
rect 12404 -3752 12415 -3699
rect 12469 -3752 12480 -3699
rect 12404 -3765 12480 -3752
rect 13472 -3714 13586 -3692
rect 8539 -3797 8643 -3783
rect 13472 -3774 13507 -3714
rect 13570 -3774 13586 -3714
rect 17250 -3699 17326 -2072
rect 19432 -2702 19544 -2697
rect 19432 -2758 19458 -2702
rect 19521 -2758 19544 -2702
rect 19432 -2761 19544 -2758
rect 18558 -2812 18642 -2798
rect 18315 -2835 18440 -2828
rect 18315 -2891 18340 -2835
rect 18412 -2891 18440 -2835
rect 18558 -2870 18570 -2812
rect 18629 -2870 18642 -2812
rect 18558 -2878 18642 -2870
rect 18315 -2905 18440 -2891
rect 17250 -3752 17261 -3699
rect 17315 -3752 17326 -3699
rect 17250 -3765 17326 -3752
rect 18233 -3716 18335 -3695
rect 13472 -3803 13586 -3774
rect 18233 -3777 18259 -3716
rect 18323 -3777 18335 -3716
rect 22096 -3699 22172 -2072
rect 24248 -2699 24360 -2697
rect 24248 -2756 24269 -2699
rect 24334 -2756 24360 -2699
rect 24248 -2761 24360 -2756
rect 23402 -2813 23491 -2796
rect 23156 -2834 23280 -2828
rect 23156 -2890 23186 -2834
rect 23258 -2890 23280 -2834
rect 23402 -2870 23416 -2813
rect 23475 -2870 23491 -2813
rect 23402 -2883 23491 -2870
rect 23156 -2905 23280 -2890
rect 26942 -3699 27018 -2072
rect 29120 -2702 29232 -2697
rect 29120 -2758 29145 -2702
rect 29206 -2758 29232 -2702
rect 29120 -2761 29232 -2758
rect 28246 -2810 28340 -2801
rect 28010 -2834 28127 -2828
rect 28010 -2890 28032 -2834
rect 28104 -2890 28127 -2834
rect 28246 -2868 28265 -2810
rect 28322 -2868 28340 -2810
rect 28246 -2881 28340 -2868
rect 28010 -2905 28127 -2890
rect 22096 -3752 22107 -3699
rect 22161 -3752 22172 -3699
rect 22096 -3765 22172 -3752
rect 23155 -3718 23270 -3699
rect 18233 -3801 18335 -3777
rect 23155 -3774 23194 -3718
rect 23253 -3774 23270 -3718
rect 26942 -3752 26953 -3699
rect 27007 -3752 27018 -3699
rect 26942 -3765 27018 -3752
rect 27965 -3714 28068 -3696
rect 23155 -3796 23270 -3774
rect 27965 -3772 27990 -3714
rect 28052 -3772 28068 -3714
rect 31788 -3699 31864 -2072
rect 33963 -2701 34077 -2697
rect 33963 -2757 33989 -2701
rect 34051 -2757 34077 -2701
rect 33963 -2761 34077 -2757
rect 33092 -2813 33180 -2801
rect 32851 -2832 32982 -2828
rect 32851 -2889 32878 -2832
rect 32950 -2889 32982 -2832
rect 33092 -2869 33110 -2813
rect 33166 -2869 33180 -2813
rect 33092 -2880 33180 -2869
rect 32851 -2905 32982 -2889
rect 31788 -3752 31799 -3699
rect 31853 -3752 31864 -3699
rect 31788 -3765 31864 -3752
rect 32843 -3714 32940 -3695
rect 27965 -3796 28068 -3772
rect 32843 -3774 32869 -3714
rect 32932 -3774 32940 -3714
rect 36634 -3699 36710 -2072
rect 38808 -2702 38920 -2697
rect 38808 -2758 38833 -2702
rect 38894 -2758 38920 -2702
rect 38808 -2761 38920 -2758
rect 37693 -2834 37824 -2828
rect 37693 -2892 37724 -2834
rect 37796 -2892 37824 -2834
rect 37693 -2905 37824 -2892
rect 36634 -3752 36645 -3699
rect 36699 -3752 36710 -3699
rect 36634 -3765 36710 -3752
rect 41480 -3699 41556 -2072
rect 41480 -3752 41491 -3699
rect 41545 -3752 41556 -3699
rect 41480 -3765 41556 -3752
rect 32843 -3788 32940 -3774
rect 7591 -3850 8083 -3839
rect 7591 -3851 8019 -3850
rect 7591 -3904 7602 -3851
rect 7656 -3903 8019 -3851
rect 8073 -3903 8083 -3850
rect 7656 -3904 8083 -3903
rect 7591 -3915 8083 -3904
rect 12437 -3850 12929 -3839
rect 12437 -3851 12865 -3850
rect 12437 -3904 12448 -3851
rect 12502 -3903 12865 -3851
rect 12919 -3903 12929 -3850
rect 12502 -3904 12929 -3903
rect 12437 -3915 12929 -3904
rect 17283 -3850 17775 -3839
rect 17283 -3851 17711 -3850
rect 17283 -3904 17294 -3851
rect 17348 -3903 17711 -3851
rect 17765 -3903 17775 -3850
rect 17348 -3904 17775 -3903
rect 17283 -3915 17775 -3904
rect 22129 -3850 22621 -3839
rect 22129 -3851 22557 -3850
rect 22129 -3904 22140 -3851
rect 22194 -3903 22557 -3851
rect 22611 -3903 22621 -3850
rect 22194 -3904 22621 -3903
rect 22129 -3915 22621 -3904
rect 26975 -3850 27467 -3839
rect 26975 -3851 27403 -3850
rect 26975 -3904 26986 -3851
rect 27040 -3903 27403 -3851
rect 27457 -3903 27467 -3850
rect 27040 -3904 27467 -3903
rect 26975 -3915 27467 -3904
rect 31821 -3850 32313 -3839
rect 31821 -3851 32249 -3850
rect 31821 -3904 31832 -3851
rect 31886 -3903 32249 -3851
rect 32303 -3903 32313 -3850
rect 31886 -3904 32313 -3903
rect 31821 -3915 32313 -3904
rect 36667 -3850 37159 -3839
rect 36667 -3851 37095 -3850
rect 36667 -3904 36678 -3851
rect 36732 -3903 37095 -3851
rect 37149 -3903 37159 -3850
rect 36732 -3904 37159 -3903
rect 36667 -3915 37159 -3904
rect 41513 -3850 42005 -3839
rect 41513 -3851 41941 -3850
rect 41513 -3904 41524 -3851
rect 41578 -3903 41941 -3851
rect 41995 -3903 42005 -3850
rect 41578 -3904 42005 -3903
rect 41513 -3915 42005 -3904
rect 7798 -4256 7874 -3915
rect 12644 -4256 12720 -3915
rect 17490 -4256 17566 -3915
rect 22336 -4256 22412 -3915
rect 27182 -4256 27258 -3915
rect 32028 -4256 32104 -3915
rect 36874 -4256 36950 -3915
rect 41720 -4256 41796 -3915
rect 7392 -4424 42616 -4256
rect 42784 -4424 42857 -4256
rect 43064 -4704 43400 -2072
rect 7504 -4872 43400 -4704
rect 4872 -5499 4984 -5497
rect 4872 -5555 4893 -5499
rect 4956 -5555 4984 -5499
rect 4872 -5561 4984 -5555
rect 4015 -5612 4108 -5609
rect 3772 -5637 3900 -5629
rect 3772 -5693 3802 -5637
rect 3874 -5693 3900 -5637
rect 4015 -5668 4035 -5612
rect 4091 -5668 4108 -5612
rect 4015 -5675 4108 -5668
rect 3772 -5705 3900 -5693
rect 3068 -5826 3150 -5773
rect 3068 -5840 3076 -5826
rect 2734 -5907 3076 -5840
rect 3146 -5907 3150 -5826
rect 2734 -5925 3150 -5907
rect 2734 -6277 2819 -5925
rect 2734 -6330 2750 -6277
rect 2740 -6351 2750 -6330
rect 2803 -6330 2819 -6277
rect 2803 -6351 2812 -6330
rect 2740 -6370 2812 -6351
rect 3077 -6512 3154 -6502
rect 3077 -6569 3087 -6512
rect 3146 -6569 3154 -6512
rect 3077 -6581 3154 -6569
rect 3660 -6507 3762 -6493
rect 3660 -6583 3691 -6507
rect 3750 -6583 3762 -6507
rect 7558 -6499 7634 -4872
rect 9744 -5498 9856 -5497
rect 9744 -5554 9772 -5498
rect 9834 -5554 9856 -5498
rect 9744 -5561 9856 -5554
rect 8860 -5613 8955 -5608
rect 8624 -5632 8757 -5627
rect 8624 -5690 8648 -5632
rect 8720 -5690 8757 -5632
rect 8860 -5670 8878 -5613
rect 8937 -5670 8955 -5613
rect 8860 -5674 8955 -5670
rect 8624 -5705 8757 -5690
rect 7558 -6552 7569 -6499
rect 7623 -6552 7634 -6499
rect 7558 -6565 7634 -6552
rect 8529 -6507 8634 -6496
rect 3660 -6600 3762 -6583
rect 8529 -6583 8565 -6507
rect 8624 -6583 8634 -6507
rect 12404 -6499 12480 -4872
rect 14560 -5501 14672 -5497
rect 14560 -5557 14580 -5501
rect 14645 -5557 14672 -5501
rect 14560 -5561 14672 -5557
rect 13701 -5613 13802 -5602
rect 13470 -5635 13601 -5627
rect 13470 -5692 13494 -5635
rect 13566 -5692 13601 -5635
rect 13701 -5669 13725 -5613
rect 13783 -5669 13802 -5613
rect 13701 -5679 13802 -5669
rect 13470 -5705 13601 -5692
rect 12404 -6552 12415 -6499
rect 12469 -6552 12480 -6499
rect 12404 -6565 12480 -6552
rect 13470 -6513 13579 -6495
rect 8529 -6597 8634 -6583
rect 13470 -6573 13506 -6513
rect 13569 -6573 13579 -6513
rect 17250 -6499 17326 -4872
rect 19432 -5502 19544 -5497
rect 19432 -5558 19458 -5502
rect 19521 -5558 19544 -5502
rect 19432 -5561 19544 -5558
rect 18556 -5607 18645 -5598
rect 18312 -5634 18442 -5627
rect 18312 -5691 18340 -5634
rect 18412 -5691 18442 -5634
rect 18556 -5671 18569 -5607
rect 18634 -5671 18645 -5607
rect 18556 -5682 18645 -5671
rect 18312 -5705 18442 -5691
rect 17250 -6552 17261 -6499
rect 17315 -6552 17326 -6499
rect 17250 -6565 17326 -6552
rect 18230 -6517 18333 -6492
rect 13470 -6597 13579 -6573
rect 18230 -6577 18253 -6517
rect 18318 -6577 18333 -6517
rect 22096 -6499 22172 -4872
rect 24248 -5499 24360 -5497
rect 24248 -5556 24269 -5499
rect 24334 -5556 24360 -5499
rect 24248 -5561 24360 -5556
rect 23404 -5610 23490 -5601
rect 23162 -5634 23290 -5627
rect 23162 -5691 23186 -5634
rect 23258 -5691 23290 -5634
rect 23404 -5671 23416 -5610
rect 23478 -5671 23490 -5610
rect 23404 -5683 23490 -5671
rect 23162 -5705 23290 -5691
rect 22096 -6552 22107 -6499
rect 22161 -6552 22172 -6499
rect 22096 -6565 22172 -6552
rect 23153 -6516 23268 -6495
rect 18230 -6599 18333 -6577
rect 23153 -6572 23194 -6516
rect 23252 -6572 23268 -6516
rect 26942 -6499 27018 -4872
rect 29120 -5502 29232 -5497
rect 29120 -5558 29145 -5502
rect 29206 -5558 29232 -5502
rect 29120 -5561 29232 -5558
rect 28251 -5611 28335 -5601
rect 28004 -5634 28132 -5628
rect 28004 -5691 28032 -5634
rect 28104 -5691 28132 -5634
rect 28251 -5668 28264 -5611
rect 28323 -5668 28335 -5611
rect 28251 -5683 28335 -5668
rect 28004 -5705 28132 -5691
rect 26942 -6552 26953 -6499
rect 27007 -6552 27018 -6499
rect 26942 -6565 27018 -6552
rect 27963 -6515 28073 -6494
rect 23153 -6597 23268 -6572
rect 27963 -6576 27985 -6515
rect 28045 -6576 28073 -6515
rect 31788 -6499 31864 -4872
rect 33963 -5501 34077 -5497
rect 33963 -5557 33989 -5501
rect 34051 -5557 34077 -5501
rect 33963 -5561 34077 -5557
rect 33096 -5611 33179 -5606
rect 32853 -5634 32974 -5627
rect 32853 -5691 32878 -5634
rect 32950 -5691 32974 -5634
rect 33096 -5669 33109 -5611
rect 33169 -5669 33179 -5611
rect 33096 -5679 33179 -5669
rect 32853 -5705 32974 -5691
rect 31788 -6552 31799 -6499
rect 31853 -6552 31864 -6499
rect 36634 -6499 36710 -4872
rect 38808 -5502 38920 -5497
rect 38808 -5558 38833 -5502
rect 38894 -5558 38920 -5502
rect 38808 -5561 38920 -5558
rect 37944 -5612 38026 -5602
rect 37944 -5668 37956 -5612
rect 38014 -5668 38026 -5612
rect 37944 -5678 38026 -5668
rect 31788 -6565 31864 -6552
rect 32851 -6517 32944 -6500
rect 27963 -6597 28073 -6576
rect 32851 -6573 32870 -6517
rect 32933 -6573 32944 -6517
rect 36634 -6552 36645 -6499
rect 36699 -6552 36710 -6499
rect 36634 -6565 36710 -6552
rect 41480 -6499 41556 -4872
rect 41480 -6552 41491 -6499
rect 41545 -6552 41556 -6499
rect 41480 -6565 41556 -6552
rect 32851 -6588 32944 -6573
rect 7591 -6650 8083 -6639
rect 7591 -6651 8019 -6650
rect 7591 -6704 7602 -6651
rect 7656 -6703 8019 -6651
rect 8073 -6703 8083 -6650
rect 7656 -6704 8083 -6703
rect 7591 -6715 8083 -6704
rect 12437 -6650 12929 -6639
rect 12437 -6651 12865 -6650
rect 12437 -6704 12448 -6651
rect 12502 -6703 12865 -6651
rect 12919 -6703 12929 -6650
rect 12502 -6704 12929 -6703
rect 12437 -6715 12929 -6704
rect 17283 -6650 17775 -6639
rect 17283 -6651 17711 -6650
rect 17283 -6704 17294 -6651
rect 17348 -6703 17711 -6651
rect 17765 -6703 17775 -6650
rect 17348 -6704 17775 -6703
rect 17283 -6715 17775 -6704
rect 22129 -6650 22621 -6639
rect 22129 -6651 22557 -6650
rect 22129 -6704 22140 -6651
rect 22194 -6703 22557 -6651
rect 22611 -6703 22621 -6650
rect 22194 -6704 22621 -6703
rect 22129 -6715 22621 -6704
rect 26975 -6650 27467 -6639
rect 26975 -6651 27403 -6650
rect 26975 -6704 26986 -6651
rect 27040 -6703 27403 -6651
rect 27457 -6703 27467 -6650
rect 27040 -6704 27467 -6703
rect 26975 -6715 27467 -6704
rect 31821 -6650 32313 -6639
rect 31821 -6651 32249 -6650
rect 31821 -6704 31832 -6651
rect 31886 -6703 32249 -6651
rect 32303 -6703 32313 -6650
rect 31886 -6704 32313 -6703
rect 31821 -6715 32313 -6704
rect 36667 -6650 37159 -6639
rect 36667 -6651 37095 -6650
rect 36667 -6704 36678 -6651
rect 36732 -6703 37095 -6651
rect 37149 -6703 37159 -6650
rect 36732 -6704 37159 -6703
rect 36667 -6715 37159 -6704
rect 41513 -6650 42005 -6639
rect 41513 -6651 41941 -6650
rect 41513 -6704 41524 -6651
rect 41578 -6703 41941 -6651
rect 41995 -6703 42005 -6650
rect 41578 -6704 42005 -6703
rect 41513 -6715 42005 -6704
rect 7798 -7056 7874 -6715
rect 12644 -7056 12720 -6715
rect 17490 -7056 17566 -6715
rect 22336 -7056 22412 -6715
rect 27182 -7056 27258 -6715
rect 32028 -7056 32104 -6715
rect 36874 -7056 36950 -6715
rect 41720 -7056 41796 -6715
rect 7392 -7224 42616 -7056
rect 42784 -7224 42857 -7056
rect 43064 -7504 43400 -4872
rect 7504 -7672 43400 -7504
rect 4872 -8299 4984 -8297
rect 4872 -8355 4893 -8299
rect 4956 -8355 4984 -8299
rect 4872 -8361 4984 -8355
rect 4013 -8413 4113 -8406
rect 3778 -8434 3891 -8429
rect 3778 -8493 3802 -8434
rect 3874 -8493 3891 -8434
rect 4013 -8469 4034 -8413
rect 4091 -8469 4113 -8413
rect 4013 -8478 4113 -8469
rect 3778 -8505 3891 -8493
rect 7558 -9299 7634 -7672
rect 9744 -8298 9856 -8297
rect 9744 -8354 9772 -8298
rect 9834 -8354 9856 -8298
rect 9744 -8361 9856 -8354
rect 8854 -8411 8968 -8405
rect 8625 -8435 8746 -8427
rect 8625 -8492 8648 -8435
rect 8720 -8492 8746 -8435
rect 8854 -8471 8878 -8411
rect 8942 -8471 8968 -8411
rect 8854 -8481 8968 -8471
rect 8625 -8505 8746 -8492
rect 3670 -9317 3776 -9299
rect 3670 -9373 3696 -9317
rect 3752 -9373 3776 -9317
rect 7558 -9352 7569 -9299
rect 7623 -9352 7634 -9299
rect 7558 -9365 7634 -9352
rect 8529 -9307 8645 -9296
rect 3286 -9400 3380 -9379
rect 3670 -9397 3776 -9373
rect 8529 -9383 8566 -9307
rect 8627 -9383 8645 -9307
rect 12404 -9299 12480 -7672
rect 14560 -8301 14672 -8297
rect 14560 -8357 14580 -8301
rect 14645 -8357 14672 -8301
rect 14560 -8361 14672 -8357
rect 13705 -8413 13804 -8401
rect 13468 -8433 13598 -8427
rect 13468 -8491 13494 -8433
rect 13566 -8491 13598 -8433
rect 13705 -8469 13726 -8413
rect 13782 -8469 13804 -8413
rect 13705 -8478 13804 -8469
rect 13468 -8505 13598 -8491
rect 12404 -9352 12415 -9299
rect 12469 -9352 12480 -9299
rect 12404 -9365 12480 -9352
rect 13467 -9314 13579 -9296
rect 3286 -9464 3298 -9400
rect 3362 -9464 3380 -9400
rect 8529 -9402 8645 -9383
rect 13467 -9373 13505 -9314
rect 13570 -9373 13579 -9314
rect 17250 -9299 17326 -7672
rect 19432 -8302 19544 -8297
rect 19432 -8358 19458 -8302
rect 19521 -8358 19544 -8302
rect 19432 -8361 19544 -8358
rect 18550 -8412 18647 -8398
rect 18312 -8433 18445 -8427
rect 18312 -8491 18340 -8433
rect 18412 -8491 18445 -8433
rect 18312 -8505 18445 -8491
rect 18550 -8470 18571 -8412
rect 18629 -8470 18647 -8412
rect 18550 -8493 18647 -8470
rect 17250 -9352 17261 -9299
rect 17315 -9352 17326 -9299
rect 17250 -9365 17326 -9352
rect 18226 -9317 18333 -9296
rect 13467 -9399 13579 -9373
rect 18226 -9376 18252 -9317
rect 18318 -9376 18333 -9317
rect 22096 -9299 22172 -7672
rect 24248 -8299 24360 -8297
rect 24248 -8356 24269 -8299
rect 24334 -8356 24360 -8299
rect 24248 -8361 24360 -8356
rect 23405 -8406 23490 -8393
rect 23159 -8434 23292 -8427
rect 23159 -8491 23186 -8434
rect 23258 -8491 23292 -8434
rect 23405 -8471 23416 -8406
rect 23479 -8471 23490 -8406
rect 23405 -8481 23490 -8471
rect 23159 -8505 23292 -8491
rect 22096 -9352 22107 -9299
rect 22161 -9352 22172 -9299
rect 22096 -9365 22172 -9352
rect 23153 -9314 23265 -9295
rect 18226 -9396 18333 -9376
rect 23153 -9373 23194 -9314
rect 23252 -9373 23265 -9314
rect 26942 -9299 27018 -7672
rect 29120 -8302 29232 -8297
rect 29120 -8358 29145 -8302
rect 29206 -8358 29232 -8302
rect 29120 -8361 29232 -8358
rect 28247 -8411 28343 -8401
rect 28008 -8433 28137 -8427
rect 28008 -8492 28032 -8433
rect 28104 -8492 28137 -8433
rect 28247 -8469 28262 -8411
rect 28323 -8469 28343 -8411
rect 28247 -8487 28343 -8469
rect 28008 -8505 28137 -8492
rect 26942 -9352 26953 -9299
rect 27007 -9352 27018 -9299
rect 26942 -9365 27018 -9352
rect 27968 -9317 28077 -9293
rect 23153 -9397 23265 -9373
rect 27968 -9375 27993 -9317
rect 28053 -9375 28077 -9317
rect 31788 -9299 31864 -7672
rect 33963 -8301 34077 -8297
rect 33963 -8357 33989 -8301
rect 34051 -8357 34077 -8301
rect 33963 -8361 34077 -8357
rect 33093 -8413 33183 -8403
rect 32853 -8434 32980 -8427
rect 32853 -8490 32878 -8434
rect 32950 -8490 32980 -8434
rect 33093 -8471 33107 -8413
rect 33166 -8471 33183 -8413
rect 33093 -8484 33183 -8471
rect 32853 -8505 32980 -8490
rect 31788 -9352 31799 -9299
rect 31853 -9352 31864 -9299
rect 36634 -9299 36710 -7672
rect 38808 -8302 38920 -8297
rect 38808 -8358 38833 -8302
rect 38894 -8358 38920 -8302
rect 38808 -8361 38920 -8358
rect 37938 -8413 38026 -8407
rect 37938 -8469 37955 -8413
rect 38013 -8469 38026 -8413
rect 37938 -8478 38026 -8469
rect 31788 -9365 31864 -9352
rect 32853 -9316 32946 -9300
rect 27968 -9397 28077 -9375
rect 32853 -9374 32867 -9316
rect 32933 -9374 32946 -9316
rect 36634 -9352 36645 -9299
rect 36699 -9352 36710 -9299
rect 36634 -9365 36710 -9352
rect 41480 -9299 41556 -7672
rect 41480 -9352 41491 -9299
rect 41545 -9352 41556 -9299
rect 41480 -9365 41556 -9352
rect 32853 -9387 32946 -9374
rect 3286 -9477 3380 -9464
rect 7591 -9450 8083 -9439
rect 7591 -9451 8019 -9450
rect 7591 -9504 7602 -9451
rect 7656 -9503 8019 -9451
rect 8073 -9503 8083 -9450
rect 7656 -9504 8083 -9503
rect 7591 -9515 8083 -9504
rect 12437 -9450 12929 -9439
rect 12437 -9451 12865 -9450
rect 12437 -9504 12448 -9451
rect 12502 -9503 12865 -9451
rect 12919 -9503 12929 -9450
rect 12502 -9504 12929 -9503
rect 12437 -9515 12929 -9504
rect 17283 -9450 17775 -9439
rect 17283 -9451 17711 -9450
rect 17283 -9504 17294 -9451
rect 17348 -9503 17711 -9451
rect 17765 -9503 17775 -9450
rect 17348 -9504 17775 -9503
rect 17283 -9515 17775 -9504
rect 22129 -9450 22621 -9439
rect 22129 -9451 22557 -9450
rect 22129 -9504 22140 -9451
rect 22194 -9503 22557 -9451
rect 22611 -9503 22621 -9450
rect 22194 -9504 22621 -9503
rect 22129 -9515 22621 -9504
rect 26975 -9450 27467 -9439
rect 26975 -9451 27403 -9450
rect 26975 -9504 26986 -9451
rect 27040 -9503 27403 -9451
rect 27457 -9503 27467 -9450
rect 27040 -9504 27467 -9503
rect 26975 -9515 27467 -9504
rect 31821 -9450 32313 -9439
rect 31821 -9451 32249 -9450
rect 31821 -9504 31832 -9451
rect 31886 -9503 32249 -9451
rect 32303 -9503 32313 -9450
rect 31886 -9504 32313 -9503
rect 31821 -9515 32313 -9504
rect 36667 -9450 37159 -9439
rect 36667 -9451 37095 -9450
rect 36667 -9504 36678 -9451
rect 36732 -9503 37095 -9451
rect 37149 -9503 37159 -9450
rect 36732 -9504 37159 -9503
rect 36667 -9515 37159 -9504
rect 41513 -9450 42005 -9439
rect 41513 -9451 41941 -9450
rect 41513 -9504 41524 -9451
rect 41578 -9503 41941 -9451
rect 41995 -9503 42005 -9450
rect 41578 -9504 42005 -9503
rect 41513 -9515 42005 -9504
rect 7798 -9856 7874 -9515
rect 12644 -9856 12720 -9515
rect 17490 -9856 17566 -9515
rect 22336 -9856 22412 -9515
rect 27182 -9856 27258 -9515
rect 32028 -9856 32104 -9515
rect 36874 -9856 36950 -9515
rect 41720 -9856 41796 -9515
rect 7392 -10024 42616 -9856
rect 42784 -10024 42857 -9856
rect 43064 -10304 43400 -7672
rect 7504 -10472 43400 -10304
rect 4872 -11099 4984 -11097
rect 4872 -11155 4893 -11099
rect 4956 -11155 4984 -11099
rect 4872 -11161 4984 -11155
rect 4013 -11212 4108 -11207
rect 3777 -11232 3902 -11227
rect 3777 -11291 3802 -11232
rect 3874 -11291 3902 -11232
rect 4013 -11268 4035 -11212
rect 4091 -11268 4108 -11212
rect 4013 -11277 4108 -11268
rect 3777 -11305 3902 -11291
rect 3090 -11421 3161 -11374
rect 3090 -11445 3096 -11421
rect 2860 -11514 3096 -11445
rect 3157 -11514 3161 -11421
rect 2860 -11517 3161 -11514
rect 2860 -11876 2932 -11517
rect 3090 -11527 3161 -11517
rect 2860 -11959 2865 -11876
rect 2926 -11959 2932 -11876
rect 2860 -11977 2932 -11959
rect 3665 -12107 3777 -12095
rect 3181 -12155 3276 -12147
rect 3181 -12228 3197 -12155
rect 3267 -12228 3276 -12155
rect 3665 -12183 3688 -12107
rect 3758 -12183 3777 -12107
rect 7558 -12099 7634 -10472
rect 9744 -11098 9856 -11097
rect 9744 -11154 9772 -11098
rect 9834 -11154 9856 -11098
rect 9744 -11161 9856 -11154
rect 8855 -11212 8956 -11201
rect 8625 -11235 8744 -11227
rect 8625 -11291 8648 -11235
rect 8720 -11291 8744 -11235
rect 8855 -11272 8874 -11212
rect 8938 -11272 8956 -11212
rect 8855 -11284 8956 -11272
rect 8625 -11305 8744 -11291
rect 7558 -12152 7569 -12099
rect 7623 -12152 7634 -12099
rect 7558 -12165 7634 -12152
rect 8523 -12114 8641 -12093
rect 3665 -12198 3777 -12183
rect 8523 -12174 8559 -12114
rect 8617 -12174 8641 -12114
rect 12404 -12099 12480 -10472
rect 14560 -11101 14672 -11097
rect 14560 -11157 14580 -11101
rect 14645 -11157 14672 -11101
rect 14560 -11161 14672 -11157
rect 13707 -11212 13797 -11202
rect 13460 -11233 13602 -11227
rect 13460 -11293 13494 -11233
rect 13566 -11293 13602 -11233
rect 13707 -11269 13726 -11212
rect 13782 -11269 13797 -11212
rect 13707 -11284 13797 -11269
rect 13460 -11305 13602 -11293
rect 12404 -12152 12415 -12099
rect 12469 -12152 12480 -12099
rect 12404 -12165 12480 -12152
rect 13474 -12116 13574 -12096
rect 8523 -12204 8641 -12174
rect 13474 -12173 13504 -12116
rect 13564 -12173 13574 -12116
rect 17250 -12099 17326 -10472
rect 19432 -11102 19544 -11097
rect 19432 -11158 19458 -11102
rect 19521 -11158 19544 -11102
rect 19432 -11161 19544 -11158
rect 18556 -11210 18647 -11195
rect 18315 -11231 18437 -11225
rect 18315 -11291 18340 -11231
rect 18412 -11291 18437 -11231
rect 18556 -11270 18571 -11210
rect 18630 -11270 18647 -11210
rect 18556 -11284 18647 -11270
rect 18315 -11305 18437 -11291
rect 17250 -12152 17261 -12099
rect 17315 -12152 17326 -12099
rect 17250 -12165 17326 -12152
rect 18221 -12118 18325 -12094
rect 13474 -12192 13574 -12173
rect 18221 -12177 18249 -12118
rect 18313 -12177 18325 -12118
rect 22096 -12099 22172 -10472
rect 24248 -11099 24360 -11097
rect 24248 -11156 24269 -11099
rect 24334 -11156 24360 -11099
rect 24248 -11161 24360 -11156
rect 23405 -11210 23490 -11197
rect 23149 -11235 23295 -11226
rect 23149 -11293 23186 -11235
rect 23258 -11293 23295 -11235
rect 23405 -11270 23417 -11210
rect 23480 -11270 23490 -11210
rect 23405 -11283 23490 -11270
rect 23149 -11305 23295 -11293
rect 22096 -12152 22107 -12099
rect 22161 -12152 22172 -12099
rect 22096 -12165 22172 -12152
rect 23150 -12113 23268 -12095
rect 18221 -12198 18325 -12177
rect 23150 -12176 23190 -12113
rect 23255 -12176 23268 -12113
rect 26942 -12099 27018 -10472
rect 29120 -11102 29232 -11097
rect 29120 -11158 29145 -11102
rect 29206 -11158 29232 -11102
rect 29120 -11161 29232 -11158
rect 28248 -11212 28335 -11204
rect 28007 -11234 28135 -11226
rect 28007 -11291 28032 -11234
rect 28104 -11291 28135 -11234
rect 28248 -11268 28264 -11212
rect 28320 -11268 28335 -11212
rect 28248 -11278 28335 -11268
rect 28007 -11305 28135 -11291
rect 26942 -12152 26953 -12099
rect 27007 -12152 27018 -12099
rect 31788 -12099 31864 -10472
rect 33963 -11101 34077 -11097
rect 33963 -11157 33989 -11101
rect 34051 -11157 34077 -11101
rect 33963 -11161 34077 -11157
rect 33095 -11212 33179 -11203
rect 32849 -11234 32983 -11226
rect 32849 -11291 32878 -11234
rect 32950 -11291 32983 -11234
rect 33095 -11268 33111 -11212
rect 33167 -11268 33179 -11212
rect 33095 -11279 33179 -11268
rect 32849 -11305 32983 -11291
rect 26942 -12165 27018 -12152
rect 27977 -12117 28074 -12100
rect 23150 -12194 23268 -12176
rect 27977 -12175 27998 -12117
rect 28058 -12175 28074 -12117
rect 31788 -12152 31799 -12099
rect 31853 -12152 31864 -12099
rect 36634 -12099 36710 -10472
rect 38808 -11102 38920 -11097
rect 38808 -11158 38833 -11102
rect 38894 -11158 38920 -11102
rect 38808 -11161 38920 -11158
rect 37941 -11213 38024 -11203
rect 37941 -11269 37956 -11213
rect 38014 -11269 38024 -11213
rect 37941 -11279 38024 -11269
rect 31788 -12165 31864 -12152
rect 32865 -12116 32956 -12100
rect 27977 -12195 28074 -12175
rect 32865 -12173 32888 -12116
rect 32944 -12173 32956 -12116
rect 36634 -12152 36645 -12099
rect 36699 -12152 36710 -12099
rect 36634 -12165 36710 -12152
rect 41480 -12099 41556 -10472
rect 41480 -12152 41491 -12099
rect 41545 -12152 41556 -12099
rect 41480 -12165 41556 -12152
rect 32865 -12190 32956 -12173
rect 3181 -12250 3276 -12228
rect 7591 -12250 8083 -12239
rect 7591 -12251 8019 -12250
rect 7591 -12304 7602 -12251
rect 7656 -12303 8019 -12251
rect 8073 -12303 8083 -12250
rect 7656 -12304 8083 -12303
rect 7591 -12315 8083 -12304
rect 12437 -12250 12929 -12239
rect 12437 -12251 12865 -12250
rect 12437 -12304 12448 -12251
rect 12502 -12303 12865 -12251
rect 12919 -12303 12929 -12250
rect 12502 -12304 12929 -12303
rect 12437 -12315 12929 -12304
rect 17283 -12250 17775 -12239
rect 17283 -12251 17711 -12250
rect 17283 -12304 17294 -12251
rect 17348 -12303 17711 -12251
rect 17765 -12303 17775 -12250
rect 17348 -12304 17775 -12303
rect 17283 -12315 17775 -12304
rect 22129 -12250 22621 -12239
rect 22129 -12251 22557 -12250
rect 22129 -12304 22140 -12251
rect 22194 -12303 22557 -12251
rect 22611 -12303 22621 -12250
rect 22194 -12304 22621 -12303
rect 22129 -12315 22621 -12304
rect 26975 -12250 27467 -12239
rect 26975 -12251 27403 -12250
rect 26975 -12304 26986 -12251
rect 27040 -12303 27403 -12251
rect 27457 -12303 27467 -12250
rect 27040 -12304 27467 -12303
rect 26975 -12315 27467 -12304
rect 31821 -12250 32313 -12239
rect 31821 -12251 32249 -12250
rect 31821 -12304 31832 -12251
rect 31886 -12303 32249 -12251
rect 32303 -12303 32313 -12250
rect 31886 -12304 32313 -12303
rect 31821 -12315 32313 -12304
rect 36667 -12250 37159 -12239
rect 36667 -12251 37095 -12250
rect 36667 -12304 36678 -12251
rect 36732 -12303 37095 -12251
rect 37149 -12303 37159 -12250
rect 36732 -12304 37159 -12303
rect 36667 -12315 37159 -12304
rect 41513 -12250 42005 -12239
rect 41513 -12251 41941 -12250
rect 41513 -12304 41524 -12251
rect 41578 -12303 41941 -12251
rect 41995 -12303 42005 -12250
rect 41578 -12304 42005 -12303
rect 41513 -12315 42005 -12304
rect 7798 -12656 7874 -12315
rect 12644 -12656 12720 -12315
rect 17490 -12656 17566 -12315
rect 22336 -12656 22412 -12315
rect 27182 -12656 27258 -12315
rect 32028 -12656 32104 -12315
rect 36874 -12656 36950 -12315
rect 41720 -12656 41796 -12315
rect 7392 -12824 42616 -12656
rect 42784 -12824 42857 -12656
rect 43064 -13104 43400 -10472
rect 7504 -13272 43400 -13104
rect 4872 -13899 4984 -13897
rect 4872 -13955 4893 -13899
rect 4956 -13955 4984 -13899
rect 4872 -13961 4984 -13955
rect 4015 -14013 4108 -14001
rect 3766 -14035 3900 -14028
rect 3766 -14091 3802 -14035
rect 3874 -14091 3900 -14035
rect 4015 -14070 4035 -14013
rect 4092 -14070 4108 -14013
rect 4015 -14078 4108 -14070
rect 3766 -14105 3900 -14091
rect 3167 -14903 3269 -14893
rect 3167 -14978 3181 -14903
rect 3257 -14978 3269 -14903
rect 3167 -15000 3269 -14978
rect 3656 -14907 3771 -14898
rect 3656 -14983 3681 -14907
rect 3746 -14983 3771 -14907
rect 7558 -14899 7634 -13272
rect 9744 -13898 9856 -13897
rect 9744 -13954 9772 -13898
rect 9834 -13954 9856 -13898
rect 9744 -13961 9856 -13954
rect 8850 -14011 8968 -13998
rect 8629 -14035 8743 -14028
rect 8629 -14091 8648 -14035
rect 8720 -14091 8743 -14035
rect 8850 -14069 8879 -14011
rect 8939 -14069 8968 -14011
rect 8850 -14080 8968 -14069
rect 8629 -14105 8743 -14091
rect 7558 -14952 7569 -14899
rect 7623 -14952 7634 -14899
rect 7558 -14965 7634 -14952
rect 8539 -14917 8649 -14896
rect 3656 -14995 3771 -14983
rect 8539 -14973 8578 -14917
rect 8636 -14973 8649 -14917
rect 12404 -14899 12480 -13272
rect 14560 -13901 14672 -13897
rect 14560 -13957 14580 -13901
rect 14645 -13957 14672 -13901
rect 14560 -13961 14672 -13957
rect 13707 -14012 13799 -14005
rect 13476 -14035 13592 -14029
rect 13476 -14092 13494 -14035
rect 13566 -14092 13592 -14035
rect 13707 -14069 13725 -14012
rect 13784 -14069 13799 -14012
rect 13707 -14079 13799 -14069
rect 13476 -14105 13592 -14092
rect 12404 -14952 12415 -14899
rect 12469 -14952 12480 -14899
rect 12404 -14965 12480 -14952
rect 13474 -14916 13578 -14897
rect 8539 -14997 8649 -14973
rect 13474 -14973 13509 -14916
rect 13568 -14973 13578 -14916
rect 17250 -14899 17326 -13272
rect 19432 -13902 19544 -13897
rect 19432 -13958 19458 -13902
rect 19521 -13958 19544 -13902
rect 19432 -13961 19544 -13958
rect 18551 -14011 18649 -13996
rect 18313 -14033 18437 -14028
rect 18313 -14090 18340 -14033
rect 18412 -14090 18437 -14033
rect 18551 -14068 18572 -14011
rect 18630 -14068 18649 -14011
rect 18551 -14088 18649 -14068
rect 18313 -14105 18437 -14090
rect 17250 -14952 17261 -14899
rect 17315 -14952 17326 -14899
rect 17250 -14965 17326 -14952
rect 18227 -14917 18340 -14891
rect 13474 -14991 13578 -14973
rect 18227 -14979 18252 -14917
rect 18316 -14979 18340 -14917
rect 22096 -14899 22172 -13272
rect 24248 -13899 24360 -13897
rect 24248 -13956 24269 -13899
rect 24334 -13956 24360 -13899
rect 24248 -13961 24360 -13956
rect 23405 -14013 23488 -14001
rect 23166 -14036 23285 -14029
rect 23166 -14092 23186 -14036
rect 23258 -14092 23285 -14036
rect 23405 -14070 23417 -14013
rect 23477 -14070 23488 -14013
rect 23405 -14080 23488 -14070
rect 23166 -14105 23285 -14092
rect 22096 -14952 22107 -14899
rect 22161 -14952 22172 -14899
rect 22096 -14965 22172 -14952
rect 23147 -14909 23265 -14892
rect 3177 -15030 3259 -15000
rect 18227 -15005 18340 -14979
rect 23147 -14974 23191 -14909
rect 23254 -14974 23265 -14909
rect 26942 -14899 27018 -13272
rect 29120 -13902 29232 -13897
rect 29120 -13958 29145 -13902
rect 29206 -13958 29232 -13902
rect 29120 -13961 29232 -13958
rect 28250 -14012 28333 -14003
rect 28008 -14037 28129 -14029
rect 28008 -14093 28032 -14037
rect 28104 -14093 28129 -14037
rect 28250 -14068 28263 -14012
rect 28321 -14068 28333 -14012
rect 28250 -14076 28333 -14068
rect 28008 -14105 28129 -14093
rect 31788 -14899 31864 -13272
rect 33963 -13901 34077 -13897
rect 33963 -13957 33989 -13901
rect 34051 -13957 34077 -13901
rect 33963 -13961 34077 -13957
rect 33095 -14012 33178 -14005
rect 32856 -14037 32973 -14029
rect 32856 -14093 32878 -14037
rect 32950 -14093 32973 -14037
rect 33095 -14069 33110 -14012
rect 33166 -14069 33178 -14012
rect 33095 -14078 33178 -14069
rect 32856 -14105 32973 -14093
rect 26942 -14952 26953 -14899
rect 27007 -14952 27018 -14899
rect 26942 -14965 27018 -14952
rect 27979 -14916 28076 -14899
rect 23147 -14996 23265 -14974
rect 27979 -14972 27997 -14916
rect 28062 -14972 28076 -14916
rect 31788 -14952 31799 -14899
rect 31853 -14952 31864 -14899
rect 36634 -14899 36710 -13272
rect 38808 -13902 38920 -13897
rect 38808 -13958 38833 -13902
rect 38894 -13958 38920 -13902
rect 38808 -13961 38920 -13958
rect 37941 -14012 38025 -14002
rect 37941 -14068 37953 -14012
rect 38013 -14068 38025 -14012
rect 37941 -14078 38025 -14068
rect 31788 -14965 31864 -14952
rect 32845 -14916 32949 -14904
rect 27979 -14989 28076 -14972
rect 32845 -14974 32866 -14916
rect 32938 -14974 32949 -14916
rect 36634 -14952 36645 -14899
rect 36699 -14952 36710 -14899
rect 36634 -14965 36710 -14952
rect 41480 -14899 41556 -13272
rect 41480 -14952 41491 -14899
rect 41545 -14952 41556 -14899
rect 41480 -14965 41556 -14952
rect 32845 -14989 32949 -14974
rect 7591 -15050 8083 -15039
rect 7591 -15051 8019 -15050
rect 7591 -15104 7602 -15051
rect 7656 -15103 8019 -15051
rect 8073 -15103 8083 -15050
rect 7656 -15104 8083 -15103
rect 7591 -15115 8083 -15104
rect 12437 -15050 12929 -15039
rect 12437 -15051 12865 -15050
rect 12437 -15104 12448 -15051
rect 12502 -15103 12865 -15051
rect 12919 -15103 12929 -15050
rect 12502 -15104 12929 -15103
rect 12437 -15115 12929 -15104
rect 17283 -15050 17775 -15039
rect 17283 -15051 17711 -15050
rect 17283 -15104 17294 -15051
rect 17348 -15103 17711 -15051
rect 17765 -15103 17775 -15050
rect 17348 -15104 17775 -15103
rect 17283 -15115 17775 -15104
rect 22129 -15050 22621 -15039
rect 22129 -15051 22557 -15050
rect 22129 -15104 22140 -15051
rect 22194 -15103 22557 -15051
rect 22611 -15103 22621 -15050
rect 22194 -15104 22621 -15103
rect 22129 -15115 22621 -15104
rect 26975 -15050 27467 -15039
rect 26975 -15051 27403 -15050
rect 26975 -15104 26986 -15051
rect 27040 -15103 27403 -15051
rect 27457 -15103 27467 -15050
rect 27040 -15104 27467 -15103
rect 26975 -15115 27467 -15104
rect 31821 -15050 32313 -15039
rect 31821 -15051 32249 -15050
rect 31821 -15104 31832 -15051
rect 31886 -15103 32249 -15051
rect 32303 -15103 32313 -15050
rect 31886 -15104 32313 -15103
rect 31821 -15115 32313 -15104
rect 36667 -15050 37159 -15039
rect 36667 -15051 37095 -15050
rect 36667 -15104 36678 -15051
rect 36732 -15103 37095 -15051
rect 37149 -15103 37159 -15050
rect 36732 -15104 37159 -15103
rect 36667 -15115 37159 -15104
rect 41513 -15050 42005 -15039
rect 41513 -15051 41941 -15050
rect 41513 -15104 41524 -15051
rect 41578 -15103 41941 -15051
rect 41995 -15103 42005 -15050
rect 41578 -15104 42005 -15103
rect 41513 -15115 42005 -15104
rect 7798 -15456 7874 -15115
rect 12644 -15456 12720 -15115
rect 17490 -15456 17566 -15115
rect 22336 -15456 22412 -15115
rect 27182 -15456 27258 -15115
rect 32028 -15456 32104 -15115
rect 36874 -15456 36950 -15115
rect 41720 -15456 41796 -15115
rect 7392 -15624 42616 -15456
rect 42784 -15624 42857 -15456
rect 43064 -15904 43400 -13272
rect 7504 -16072 43400 -15904
rect 4872 -16699 4984 -16697
rect 4872 -16755 4893 -16699
rect 4956 -16755 4984 -16699
rect 4872 -16761 4984 -16755
rect 3174 -16806 3256 -16779
rect 3174 -16883 3181 -16806
rect 3251 -16883 3256 -16806
rect 4018 -16812 4107 -16806
rect 3174 -16910 3256 -16883
rect 3779 -16835 3900 -16829
rect 3779 -16891 3802 -16835
rect 3874 -16891 3900 -16835
rect 4018 -16868 4034 -16812
rect 4090 -16868 4107 -16812
rect 4018 -16876 4107 -16868
rect 3779 -16905 3900 -16891
rect 3180 -17099 3252 -16910
rect 2844 -17171 3256 -17099
rect 2844 -17716 2916 -17171
rect 2844 -17778 2850 -17716
rect 2911 -17778 2916 -17716
rect 2844 -17790 2916 -17778
rect 3664 -17707 3776 -17696
rect 3664 -17783 3692 -17707
rect 3760 -17783 3776 -17707
rect 7558 -17699 7634 -16072
rect 9744 -16698 9856 -16697
rect 9744 -16754 9772 -16698
rect 9834 -16754 9856 -16698
rect 9744 -16761 9856 -16754
rect 8857 -16812 8959 -16805
rect 8626 -16836 8745 -16828
rect 8626 -16892 8648 -16836
rect 8720 -16892 8745 -16836
rect 8857 -16870 8879 -16812
rect 8938 -16870 8959 -16812
rect 8857 -16879 8959 -16870
rect 8626 -16905 8745 -16892
rect 7558 -17752 7569 -17699
rect 7623 -17752 7634 -17699
rect 7558 -17765 7634 -17752
rect 8538 -17717 8646 -17693
rect 3664 -17796 3776 -17783
rect 8538 -17775 8570 -17717
rect 8630 -17775 8646 -17717
rect 12404 -17699 12480 -16072
rect 14560 -16701 14672 -16697
rect 14560 -16757 14580 -16701
rect 14645 -16757 14672 -16701
rect 14560 -16761 14672 -16757
rect 13710 -16812 13795 -16806
rect 13473 -16835 13589 -16829
rect 13473 -16891 13494 -16835
rect 13566 -16891 13589 -16835
rect 13710 -16869 13726 -16812
rect 13785 -16869 13795 -16812
rect 13710 -16881 13795 -16869
rect 13473 -16905 13589 -16891
rect 17250 -17699 17326 -16072
rect 19432 -16702 19544 -16697
rect 19432 -16758 19458 -16702
rect 19521 -16758 19544 -16702
rect 19432 -16761 19544 -16758
rect 18558 -16810 18643 -16799
rect 18321 -16836 18434 -16828
rect 18321 -16892 18340 -16836
rect 18412 -16892 18434 -16836
rect 18558 -16869 18572 -16810
rect 18630 -16869 18643 -16810
rect 18558 -16884 18643 -16869
rect 18321 -16905 18434 -16892
rect 12404 -17752 12415 -17699
rect 12469 -17752 12480 -17699
rect 12404 -17765 12480 -17752
rect 13483 -17715 13572 -17699
rect 8538 -17798 8646 -17775
rect 13483 -17771 13505 -17715
rect 13561 -17771 13572 -17715
rect 17250 -17752 17261 -17699
rect 17315 -17752 17326 -17699
rect 17250 -17765 17326 -17752
rect 18221 -17715 18335 -17695
rect 13483 -17793 13572 -17771
rect 18221 -17776 18250 -17715
rect 18318 -17776 18335 -17715
rect 22096 -17699 22172 -16072
rect 24248 -16699 24360 -16697
rect 24248 -16756 24269 -16699
rect 24334 -16756 24360 -16699
rect 24248 -16761 24360 -16756
rect 23406 -16811 23491 -16801
rect 23168 -16837 23286 -16829
rect 23168 -16893 23186 -16837
rect 23258 -16893 23286 -16837
rect 23406 -16870 23415 -16811
rect 23478 -16870 23491 -16811
rect 23406 -16880 23491 -16870
rect 23168 -16905 23286 -16893
rect 22096 -17752 22107 -17699
rect 22161 -17752 22172 -17699
rect 22096 -17765 22172 -17752
rect 23153 -17712 23267 -17694
rect 18221 -17796 18335 -17776
rect 23153 -17778 23191 -17712
rect 23251 -17778 23267 -17712
rect 26942 -17699 27018 -16072
rect 29120 -16702 29232 -16697
rect 29120 -16758 29145 -16702
rect 29206 -16758 29232 -16702
rect 29120 -16761 29232 -16758
rect 28249 -16811 28334 -16804
rect 28013 -16837 28131 -16829
rect 28013 -16893 28032 -16837
rect 28104 -16893 28131 -16837
rect 28249 -16867 28265 -16811
rect 28323 -16867 28334 -16811
rect 28249 -16875 28334 -16867
rect 28013 -16905 28131 -16893
rect 26942 -17752 26953 -17699
rect 27007 -17752 27018 -17699
rect 26942 -17765 27018 -17752
rect 27983 -17712 28077 -17698
rect 23153 -17798 23267 -17778
rect 27983 -17769 27999 -17712
rect 28060 -17769 28077 -17712
rect 31788 -17699 31864 -16072
rect 33963 -16701 34077 -16697
rect 33963 -16757 33989 -16701
rect 34051 -16757 34077 -16701
rect 33963 -16761 34077 -16757
rect 33096 -16813 33184 -16801
rect 32857 -16835 32983 -16829
rect 32857 -16893 32878 -16835
rect 32950 -16893 32983 -16835
rect 33096 -16870 33109 -16813
rect 33167 -16870 33184 -16813
rect 33096 -16878 33184 -16870
rect 32857 -16905 32983 -16893
rect 31788 -17752 31799 -17699
rect 31853 -17752 31864 -17699
rect 36634 -17699 36710 -16072
rect 38808 -16702 38920 -16697
rect 38808 -16758 38833 -16702
rect 38894 -16758 38920 -16702
rect 38808 -16761 38920 -16758
rect 37943 -16808 38025 -16798
rect 37943 -16870 37953 -16808
rect 38015 -16870 38025 -16808
rect 37943 -16880 38025 -16870
rect 31788 -17765 31864 -17752
rect 32850 -17715 32945 -17702
rect 27983 -17787 28077 -17769
rect 32850 -17775 32868 -17715
rect 32935 -17775 32945 -17715
rect 36634 -17752 36645 -17699
rect 36699 -17752 36710 -17699
rect 36634 -17765 36710 -17752
rect 41480 -17699 41556 -16072
rect 41480 -17752 41491 -17699
rect 41545 -17752 41556 -17699
rect 41480 -17765 41556 -17752
rect 32850 -17791 32945 -17775
rect 7591 -17850 8083 -17839
rect 7591 -17851 8019 -17850
rect 7591 -17904 7602 -17851
rect 7656 -17903 8019 -17851
rect 8073 -17903 8083 -17850
rect 7656 -17904 8083 -17903
rect 7591 -17915 8083 -17904
rect 12437 -17850 12929 -17839
rect 12437 -17851 12865 -17850
rect 12437 -17904 12448 -17851
rect 12502 -17903 12865 -17851
rect 12919 -17903 12929 -17850
rect 12502 -17904 12929 -17903
rect 12437 -17915 12929 -17904
rect 17283 -17850 17775 -17839
rect 17283 -17851 17711 -17850
rect 17283 -17904 17294 -17851
rect 17348 -17903 17711 -17851
rect 17765 -17903 17775 -17850
rect 17348 -17904 17775 -17903
rect 17283 -17915 17775 -17904
rect 22129 -17850 22621 -17839
rect 22129 -17851 22557 -17850
rect 22129 -17904 22140 -17851
rect 22194 -17903 22557 -17851
rect 22611 -17903 22621 -17850
rect 22194 -17904 22621 -17903
rect 22129 -17915 22621 -17904
rect 26975 -17850 27467 -17839
rect 26975 -17851 27403 -17850
rect 26975 -17904 26986 -17851
rect 27040 -17903 27403 -17851
rect 27457 -17903 27467 -17850
rect 27040 -17904 27467 -17903
rect 26975 -17915 27467 -17904
rect 31821 -17850 32313 -17839
rect 31821 -17851 32249 -17850
rect 31821 -17904 31832 -17851
rect 31886 -17903 32249 -17851
rect 32303 -17903 32313 -17850
rect 31886 -17904 32313 -17903
rect 31821 -17915 32313 -17904
rect 36667 -17850 37159 -17839
rect 36667 -17851 37095 -17850
rect 36667 -17904 36678 -17851
rect 36732 -17903 37095 -17851
rect 37149 -17903 37159 -17850
rect 36732 -17904 37159 -17903
rect 36667 -17915 37159 -17904
rect 41513 -17850 42005 -17839
rect 41513 -17851 41941 -17850
rect 41513 -17904 41524 -17851
rect 41578 -17903 41941 -17851
rect 41995 -17903 42005 -17850
rect 41578 -17904 42005 -17903
rect 41513 -17915 42005 -17904
rect 7798 -18256 7874 -17915
rect 12644 -18256 12720 -17915
rect 17490 -18256 17566 -17915
rect 22336 -18256 22412 -17915
rect 27182 -18256 27258 -17915
rect 32028 -18256 32104 -17915
rect 36874 -18256 36950 -17915
rect 41720 -18256 41796 -17915
rect 7392 -18424 42616 -18256
rect 42784 -18424 42857 -18256
rect 43064 -18704 43400 -16072
rect 7504 -18872 43400 -18704
rect 4872 -19499 4984 -19497
rect 4872 -19555 4893 -19499
rect 4956 -19555 4984 -19499
rect 4872 -19561 4984 -19555
rect 4018 -19613 4107 -19608
rect 4018 -19669 4034 -19613
rect 4091 -19669 4107 -19613
rect 4018 -19678 4107 -19669
rect 3664 -20507 3772 -20496
rect 3664 -20583 3696 -20507
rect 3752 -20583 3772 -20507
rect 7558 -20499 7634 -18872
rect 9744 -19498 9856 -19497
rect 9744 -19554 9772 -19498
rect 9834 -19554 9856 -19498
rect 9744 -19561 9856 -19554
rect 8862 -19612 8956 -19603
rect 8862 -19668 8881 -19612
rect 8939 -19668 8956 -19612
rect 8862 -19678 8956 -19668
rect 7558 -20552 7569 -20499
rect 7623 -20552 7634 -20499
rect 7558 -20565 7634 -20552
rect 8532 -20514 8651 -20494
rect 3664 -20596 3772 -20583
rect 8532 -20573 8563 -20514
rect 8625 -20573 8651 -20514
rect 12404 -20499 12480 -18872
rect 14560 -19501 14672 -19497
rect 14560 -19557 14580 -19501
rect 14645 -19557 14672 -19501
rect 14560 -19561 14672 -19557
rect 13713 -19612 13794 -19602
rect 13713 -19668 13727 -19612
rect 13784 -19668 13794 -19612
rect 13713 -19676 13794 -19668
rect 12404 -20552 12415 -20499
rect 12469 -20552 12480 -20499
rect 17250 -20499 17326 -18872
rect 19432 -19502 19544 -19497
rect 19432 -19558 19458 -19502
rect 19521 -19558 19544 -19502
rect 19432 -19561 19544 -19558
rect 18555 -19613 18649 -19595
rect 18555 -19669 18573 -19613
rect 18630 -19669 18649 -19613
rect 18555 -19683 18649 -19669
rect 12404 -20565 12480 -20552
rect 13484 -20515 13581 -20501
rect 8532 -20601 8651 -20573
rect 13484 -20571 13513 -20515
rect 13571 -20571 13581 -20515
rect 17250 -20552 17261 -20499
rect 17315 -20552 17326 -20499
rect 17250 -20565 17326 -20552
rect 18223 -20518 18334 -20497
rect 13484 -20589 13581 -20571
rect 18223 -20580 18251 -20518
rect 18315 -20580 18334 -20518
rect 22096 -20499 22172 -18872
rect 24248 -19499 24360 -19497
rect 24248 -19556 24269 -19499
rect 24334 -19556 24360 -19499
rect 24248 -19561 24360 -19556
rect 23404 -19612 23485 -19605
rect 23404 -19669 23417 -19612
rect 23476 -19669 23485 -19612
rect 23404 -19679 23485 -19669
rect 22096 -20552 22107 -20499
rect 22161 -20552 22172 -20499
rect 22096 -20565 22172 -20552
rect 23162 -20514 23270 -20496
rect 18223 -20598 18334 -20580
rect 23162 -20577 23193 -20514
rect 23253 -20577 23270 -20514
rect 26942 -20499 27018 -18872
rect 29120 -19502 29232 -19497
rect 29120 -19558 29145 -19502
rect 29206 -19558 29232 -19502
rect 29120 -19561 29232 -19558
rect 28246 -19612 28338 -19599
rect 28246 -19669 28262 -19612
rect 28319 -19669 28338 -19612
rect 28246 -19681 28338 -19669
rect 26942 -20552 26953 -20499
rect 27007 -20552 27018 -20499
rect 26942 -20565 27018 -20552
rect 27983 -20517 28072 -20496
rect 23162 -20597 23270 -20577
rect 27983 -20574 27998 -20517
rect 28059 -20574 28072 -20517
rect 31788 -20499 31864 -18872
rect 33963 -19501 34077 -19497
rect 33963 -19557 33989 -19501
rect 34051 -19557 34077 -19501
rect 33963 -19561 34077 -19557
rect 33090 -19611 33189 -19600
rect 33090 -19670 33108 -19611
rect 33170 -19670 33189 -19611
rect 33090 -19685 33189 -19670
rect 31788 -20552 31799 -20499
rect 31853 -20552 31864 -20499
rect 36634 -20499 36710 -18872
rect 38744 -18873 38996 -18872
rect 43064 -19219 43400 -18872
rect 31788 -20565 31864 -20552
rect 32859 -20517 32943 -20503
rect 27983 -20587 28072 -20574
rect 32859 -20574 32869 -20517
rect 32932 -20574 32943 -20517
rect 36634 -20552 36645 -20499
rect 36699 -20552 36710 -20499
rect 36634 -20565 36710 -20552
rect 32859 -20586 32943 -20574
rect 7591 -20650 8083 -20639
rect 7591 -20651 8019 -20650
rect 7591 -20704 7602 -20651
rect 7656 -20703 8019 -20651
rect 8073 -20703 8083 -20650
rect 7656 -20704 8083 -20703
rect 7591 -20715 8083 -20704
rect 12437 -20650 12929 -20639
rect 12437 -20651 12865 -20650
rect 12437 -20704 12448 -20651
rect 12502 -20703 12865 -20651
rect 12919 -20703 12929 -20650
rect 12502 -20704 12929 -20703
rect 12437 -20715 12929 -20704
rect 17283 -20650 17775 -20639
rect 17283 -20651 17711 -20650
rect 17283 -20704 17294 -20651
rect 17348 -20703 17711 -20651
rect 17765 -20703 17775 -20650
rect 17348 -20704 17775 -20703
rect 17283 -20715 17775 -20704
rect 22129 -20650 22621 -20639
rect 22129 -20651 22557 -20650
rect 22129 -20704 22140 -20651
rect 22194 -20703 22557 -20651
rect 22611 -20703 22621 -20650
rect 22194 -20704 22621 -20703
rect 22129 -20715 22621 -20704
rect 26975 -20650 27467 -20639
rect 26975 -20651 27403 -20650
rect 26975 -20704 26986 -20651
rect 27040 -20703 27403 -20651
rect 27457 -20703 27467 -20650
rect 27040 -20704 27467 -20703
rect 26975 -20715 27467 -20704
rect 31821 -20650 32313 -20639
rect 31821 -20651 32249 -20650
rect 31821 -20704 31832 -20651
rect 31886 -20703 32249 -20651
rect 32303 -20703 32313 -20650
rect 31886 -20704 32313 -20703
rect 31821 -20715 32313 -20704
rect 36667 -20650 37159 -20639
rect 36667 -20651 37095 -20650
rect 36667 -20704 36678 -20651
rect 36732 -20703 37095 -20651
rect 37149 -20703 37159 -20650
rect 36732 -20704 37159 -20703
rect 36667 -20715 37159 -20704
rect 7798 -21056 7874 -20715
rect 12644 -21056 12720 -20715
rect 17490 -21056 17566 -20715
rect 22336 -21056 22412 -20715
rect 27182 -21056 27258 -20715
rect 32028 -21056 32104 -20715
rect 36874 -21056 36950 -20715
rect 7392 -21224 42616 -21056
rect 42785 -21224 42898 -21056
<< via2 >>
rect 3696 2436 3752 2492
rect 8568 2436 8624 2492
rect 13496 2438 13552 2494
rect 18256 2435 18312 2491
rect 23184 2436 23240 2492
rect 28000 2441 28056 2497
rect 32872 2408 32928 2464
rect 13716 1273 13780 1278
rect 13716 1206 13719 1273
rect 13719 1206 13776 1273
rect 13776 1206 13780 1273
rect 13716 1203 13780 1206
rect 18562 1254 18631 1257
rect 18562 1188 18565 1254
rect 18565 1188 18626 1254
rect 18626 1188 18631 1254
rect 18562 1185 18631 1188
rect 23403 1298 23468 1301
rect 23403 1229 23407 1298
rect 23407 1229 23464 1298
rect 23464 1229 23468 1298
rect 23403 1223 23468 1229
rect 28271 1287 28344 1291
rect 28271 1224 28280 1287
rect 28280 1224 28337 1287
rect 28337 1224 28344 1287
rect 28271 1218 28344 1224
rect 33095 1202 33156 1262
rect 6718 883 6790 888
rect 6718 822 6722 883
rect 6722 822 6785 883
rect 6785 822 6790 883
rect 6718 819 6790 822
rect 4029 485 4032 537
rect 4032 485 4088 537
rect 4088 485 4093 537
rect 4029 480 4093 485
rect 3802 -93 3874 -37
rect 4033 -15 4092 -13
rect 4033 -67 4035 -15
rect 4035 -67 4089 -15
rect 4089 -67 4092 -15
rect 4033 -69 4092 -67
rect 3110 -924 3168 -922
rect 3110 -977 3112 -924
rect 3112 -977 3165 -924
rect 3165 -977 3168 -924
rect 3110 -980 3168 -977
rect 3696 -983 3700 -907
rect 3700 -983 3768 -907
rect 3768 -983 3774 -907
rect 8648 -93 8720 -36
rect 8880 -14 8938 -12
rect 8880 -66 8882 -14
rect 8882 -66 8934 -14
rect 8934 -66 8938 -14
rect 8880 -68 8938 -66
rect 8574 -983 8632 -907
rect 13494 -38 13566 -37
rect 13494 -93 13566 -38
rect 13725 -15 13784 -13
rect 13725 -67 13727 -15
rect 13727 -67 13782 -15
rect 13782 -67 13784 -15
rect 13725 -69 13784 -67
rect 13505 -974 13567 -916
rect 18340 -90 18412 -34
rect 18570 -15 18632 -12
rect 18570 -68 18573 -15
rect 18573 -68 18628 -15
rect 18628 -68 18632 -15
rect 18570 -70 18632 -68
rect 18256 -918 18315 -915
rect 18256 -970 18259 -918
rect 18259 -970 18311 -918
rect 18311 -970 18315 -918
rect 18256 -972 18315 -970
rect 23186 -33 23258 -32
rect 23186 -88 23258 -33
rect 23418 -14 23476 -12
rect 23418 -67 23420 -14
rect 23420 -67 23474 -14
rect 23474 -67 23476 -14
rect 23418 -69 23476 -67
rect 23194 -916 23260 -913
rect 23194 -968 23199 -916
rect 23199 -968 23256 -916
rect 23256 -968 23260 -916
rect 23194 -971 23260 -968
rect 28032 -34 28104 -33
rect 28032 -89 28104 -34
rect 28262 -15 28325 -13
rect 28262 -67 28264 -15
rect 28264 -67 28322 -15
rect 28322 -67 28325 -15
rect 28262 -69 28325 -67
rect 27999 -918 28058 -915
rect 27999 -971 28001 -918
rect 28001 -971 28056 -918
rect 28056 -971 28058 -918
rect 27999 -975 28058 -971
rect 32878 -91 32950 -35
rect 33109 -15 33168 -13
rect 33109 -68 33111 -15
rect 33111 -68 33166 -15
rect 33166 -68 33168 -15
rect 33109 -70 33168 -68
rect 32869 -972 32932 -915
rect 37955 -14 38012 -13
rect 37955 -66 37959 -14
rect 37959 -66 38011 -14
rect 38011 -66 38012 -14
rect 37955 -69 38012 -66
rect 42616 -1624 42784 -1456
rect 4893 -2702 4956 -2699
rect 4893 -2755 4956 -2702
rect 3802 -2891 3874 -2835
rect 4035 -2814 4092 -2812
rect 4035 -2867 4037 -2814
rect 4037 -2867 4090 -2814
rect 4090 -2867 4092 -2814
rect 4035 -2868 4092 -2867
rect 3092 -3721 3151 -3720
rect 3092 -3778 3095 -3721
rect 3095 -3778 3148 -3721
rect 3148 -3778 3151 -3721
rect 3092 -3780 3151 -3778
rect 3687 -3783 3755 -3707
rect 9772 -2701 9834 -2698
rect 9772 -2754 9834 -2701
rect 8648 -2893 8720 -2837
rect 8879 -2815 8938 -2812
rect 8879 -2867 8882 -2815
rect 8882 -2867 8936 -2815
rect 8936 -2867 8938 -2815
rect 8879 -2870 8938 -2867
rect 8568 -3783 8628 -3707
rect 14580 -2705 14645 -2701
rect 14580 -2757 14645 -2705
rect 13494 -2892 13566 -2835
rect 13725 -2814 13784 -2812
rect 13725 -2867 13727 -2814
rect 13727 -2867 13782 -2814
rect 13782 -2867 13784 -2814
rect 13725 -2869 13784 -2867
rect 13507 -3717 13570 -3714
rect 13507 -3772 13510 -3717
rect 13510 -3772 13566 -3717
rect 13566 -3772 13570 -3717
rect 13507 -3774 13570 -3772
rect 19458 -2706 19521 -2702
rect 19458 -2758 19521 -2706
rect 18340 -2891 18412 -2835
rect 18570 -2815 18629 -2812
rect 18570 -2867 18573 -2815
rect 18573 -2867 18627 -2815
rect 18627 -2867 18629 -2815
rect 18570 -2870 18629 -2867
rect 18259 -3719 18323 -3716
rect 18259 -3773 18261 -3719
rect 18261 -3773 18319 -3719
rect 18319 -3773 18323 -3719
rect 18259 -3777 18323 -3773
rect 24269 -2703 24334 -2699
rect 24269 -2756 24334 -2703
rect 23186 -2890 23258 -2834
rect 23416 -2815 23475 -2813
rect 23416 -2868 23418 -2815
rect 23418 -2868 23472 -2815
rect 23472 -2868 23475 -2815
rect 23416 -2870 23475 -2868
rect 29145 -2705 29206 -2702
rect 29145 -2758 29206 -2705
rect 28032 -2890 28104 -2834
rect 28265 -2812 28322 -2810
rect 28265 -2866 28267 -2812
rect 28267 -2866 28320 -2812
rect 28320 -2866 28322 -2812
rect 28265 -2868 28322 -2866
rect 23194 -3774 23253 -3718
rect 27990 -3718 28052 -3714
rect 27990 -3770 27993 -3718
rect 27993 -3770 28049 -3718
rect 28049 -3770 28052 -3718
rect 27990 -3772 28052 -3770
rect 33989 -2705 34051 -2701
rect 33989 -2757 34051 -2705
rect 32878 -2889 32950 -2832
rect 33110 -2815 33166 -2813
rect 33110 -2867 33112 -2815
rect 33112 -2867 33164 -2815
rect 33164 -2867 33166 -2815
rect 33110 -2869 33166 -2867
rect 32869 -3774 32932 -3714
rect 38833 -2706 38894 -2702
rect 38833 -2758 38894 -2706
rect 37724 -2892 37796 -2834
rect 42616 -4424 42784 -4256
rect 4893 -5502 4956 -5499
rect 4893 -5555 4956 -5502
rect 3802 -5693 3874 -5637
rect 4035 -5614 4091 -5612
rect 4035 -5666 4037 -5614
rect 4037 -5666 4089 -5614
rect 4089 -5666 4091 -5614
rect 4035 -5668 4091 -5666
rect 3087 -6514 3146 -6512
rect 3087 -6566 3091 -6514
rect 3091 -6566 3143 -6514
rect 3143 -6566 3146 -6514
rect 3087 -6569 3146 -6566
rect 3691 -6583 3750 -6507
rect 9772 -5501 9834 -5498
rect 9772 -5554 9834 -5501
rect 8648 -5690 8720 -5632
rect 8878 -5615 8937 -5613
rect 8878 -5667 8882 -5615
rect 8882 -5667 8935 -5615
rect 8935 -5667 8937 -5615
rect 8878 -5670 8937 -5667
rect 8565 -6583 8624 -6507
rect 14580 -5505 14645 -5501
rect 14580 -5557 14645 -5505
rect 13494 -5692 13566 -5635
rect 13725 -5615 13783 -5613
rect 13725 -5667 13728 -5615
rect 13728 -5667 13780 -5615
rect 13780 -5667 13783 -5615
rect 13725 -5669 13783 -5667
rect 13506 -6515 13569 -6513
rect 13506 -6571 13508 -6515
rect 13508 -6571 13566 -6515
rect 13566 -6571 13569 -6515
rect 13506 -6573 13569 -6571
rect 19458 -5506 19521 -5502
rect 19458 -5558 19521 -5506
rect 18340 -5691 18412 -5634
rect 18569 -5612 18634 -5607
rect 18569 -5667 18574 -5612
rect 18574 -5667 18629 -5612
rect 18629 -5667 18634 -5612
rect 18569 -5671 18634 -5667
rect 18253 -6520 18318 -6517
rect 18253 -6573 18257 -6520
rect 18257 -6573 18315 -6520
rect 18315 -6573 18318 -6520
rect 18253 -6577 18318 -6573
rect 24269 -5503 24334 -5499
rect 24269 -5556 24334 -5503
rect 23186 -5691 23258 -5634
rect 23416 -5614 23478 -5610
rect 23416 -5667 23420 -5614
rect 23420 -5667 23473 -5614
rect 23473 -5667 23478 -5614
rect 23416 -5671 23478 -5667
rect 23194 -6517 23252 -6516
rect 23194 -6572 23250 -6517
rect 23250 -6572 23252 -6517
rect 29145 -5505 29206 -5502
rect 29145 -5558 29206 -5505
rect 28032 -5691 28104 -5634
rect 28264 -5614 28323 -5611
rect 28264 -5666 28267 -5614
rect 28267 -5666 28319 -5614
rect 28319 -5666 28323 -5614
rect 28264 -5668 28323 -5666
rect 27985 -6519 28045 -6515
rect 27985 -6574 27989 -6519
rect 27989 -6574 28042 -6519
rect 28042 -6574 28045 -6519
rect 27985 -6576 28045 -6574
rect 33989 -5505 34051 -5501
rect 33989 -5557 34051 -5505
rect 32878 -5691 32950 -5634
rect 33109 -5614 33169 -5611
rect 33109 -5667 33111 -5614
rect 33111 -5667 33165 -5614
rect 33165 -5667 33169 -5614
rect 33109 -5669 33169 -5667
rect 38833 -5506 38894 -5502
rect 38833 -5558 38894 -5506
rect 37956 -5614 38014 -5612
rect 37956 -5666 37959 -5614
rect 37959 -5666 38011 -5614
rect 38011 -5666 38014 -5614
rect 37956 -5668 38014 -5666
rect 32870 -6518 32933 -6517
rect 32870 -6573 32933 -6518
rect 42616 -7224 42784 -7056
rect 4893 -8302 4956 -8299
rect 4893 -8355 4956 -8302
rect 3802 -8493 3874 -8434
rect 4034 -8415 4091 -8413
rect 4034 -8467 4036 -8415
rect 4036 -8467 4089 -8415
rect 4089 -8467 4091 -8415
rect 4034 -8469 4091 -8467
rect 9772 -8301 9834 -8298
rect 9772 -8354 9834 -8301
rect 8648 -8492 8720 -8435
rect 8878 -8414 8942 -8411
rect 8878 -8469 8882 -8414
rect 8882 -8469 8938 -8414
rect 8938 -8469 8942 -8414
rect 8878 -8471 8942 -8469
rect 3696 -9373 3752 -9317
rect 8566 -9383 8627 -9307
rect 14580 -8305 14645 -8301
rect 14580 -8357 14645 -8305
rect 13494 -8491 13566 -8433
rect 13726 -8415 13782 -8413
rect 13726 -8467 13728 -8415
rect 13728 -8467 13780 -8415
rect 13780 -8467 13782 -8415
rect 13726 -8469 13782 -8467
rect 3298 -9464 3362 -9400
rect 13505 -9316 13570 -9314
rect 13505 -9371 13510 -9316
rect 13510 -9371 13567 -9316
rect 13567 -9371 13570 -9316
rect 13505 -9373 13570 -9371
rect 19458 -8306 19521 -8302
rect 19458 -8358 19521 -8306
rect 18340 -8491 18412 -8433
rect 18571 -8470 18629 -8412
rect 18252 -9321 18318 -9317
rect 18252 -9373 18256 -9321
rect 18256 -9373 18314 -9321
rect 18314 -9373 18318 -9321
rect 18252 -9376 18318 -9373
rect 24269 -8303 24334 -8299
rect 24269 -8356 24334 -8303
rect 23186 -8491 23258 -8434
rect 23416 -8413 23479 -8406
rect 23416 -8468 23420 -8413
rect 23420 -8468 23475 -8413
rect 23475 -8468 23479 -8413
rect 23416 -8471 23479 -8468
rect 23194 -9316 23252 -9314
rect 23194 -9371 23196 -9316
rect 23196 -9371 23250 -9316
rect 23250 -9371 23252 -9316
rect 23194 -9373 23252 -9371
rect 29145 -8305 29206 -8302
rect 29145 -8358 29206 -8305
rect 28032 -8492 28104 -8433
rect 28262 -8413 28323 -8411
rect 28262 -8467 28264 -8413
rect 28264 -8467 28321 -8413
rect 28321 -8467 28323 -8413
rect 28262 -8469 28323 -8467
rect 27993 -9375 28053 -9317
rect 33989 -8305 34051 -8301
rect 33989 -8357 34051 -8305
rect 32878 -8490 32950 -8434
rect 33107 -8414 33166 -8413
rect 33107 -8469 33110 -8414
rect 33110 -8469 33165 -8414
rect 33165 -8469 33166 -8414
rect 33107 -8471 33166 -8469
rect 38833 -8306 38894 -8302
rect 38833 -8358 38894 -8306
rect 37955 -8415 38013 -8413
rect 37955 -8467 37958 -8415
rect 37958 -8467 38010 -8415
rect 38010 -8467 38013 -8415
rect 37955 -8469 38013 -8467
rect 32867 -9317 32933 -9316
rect 32867 -9372 32868 -9317
rect 32868 -9372 32932 -9317
rect 32932 -9372 32933 -9317
rect 32867 -9374 32933 -9372
rect 42616 -10024 42784 -9856
rect 4893 -11102 4956 -11099
rect 4893 -11155 4956 -11102
rect 3802 -11291 3874 -11232
rect 4035 -11214 4091 -11212
rect 4035 -11266 4037 -11214
rect 4037 -11266 4089 -11214
rect 4089 -11266 4091 -11214
rect 4035 -11268 4091 -11266
rect 3197 -12159 3267 -12155
rect 3197 -12225 3202 -12159
rect 3202 -12225 3262 -12159
rect 3262 -12225 3267 -12159
rect 3197 -12228 3267 -12225
rect 3688 -12183 3758 -12107
rect 9772 -11101 9834 -11098
rect 9772 -11154 9834 -11101
rect 8648 -11291 8720 -11235
rect 8874 -11272 8938 -11212
rect 8559 -12118 8617 -12114
rect 8559 -12171 8562 -12118
rect 8562 -12171 8614 -12118
rect 8614 -12171 8617 -12118
rect 8559 -12174 8617 -12171
rect 14580 -11105 14645 -11101
rect 14580 -11157 14645 -11105
rect 13494 -11293 13566 -11233
rect 13726 -11214 13782 -11212
rect 13726 -11266 13728 -11214
rect 13728 -11266 13780 -11214
rect 13780 -11266 13782 -11214
rect 13726 -11269 13782 -11266
rect 13504 -12119 13564 -12116
rect 13504 -12171 13506 -12119
rect 13506 -12171 13560 -12119
rect 13560 -12171 13564 -12119
rect 13504 -12173 13564 -12171
rect 19458 -11106 19521 -11102
rect 19458 -11158 19521 -11106
rect 18340 -11291 18412 -11231
rect 18571 -11213 18630 -11210
rect 18571 -11268 18573 -11213
rect 18573 -11268 18626 -11213
rect 18626 -11268 18630 -11213
rect 18571 -11270 18630 -11268
rect 18249 -12121 18313 -12118
rect 18249 -12174 18253 -12121
rect 18253 -12174 18309 -12121
rect 18309 -12174 18313 -12121
rect 18249 -12177 18313 -12174
rect 24269 -11103 24334 -11099
rect 24269 -11156 24334 -11103
rect 23186 -11293 23258 -11235
rect 23417 -11213 23480 -11210
rect 23417 -11267 23420 -11213
rect 23420 -11267 23477 -11213
rect 23477 -11267 23480 -11213
rect 23417 -11270 23480 -11267
rect 23190 -12116 23255 -12113
rect 23190 -12173 23192 -12116
rect 23192 -12173 23252 -12116
rect 23252 -12173 23255 -12116
rect 23190 -12176 23255 -12173
rect 29145 -11105 29206 -11102
rect 29145 -11158 29206 -11105
rect 28032 -11291 28104 -11234
rect 28264 -11214 28320 -11212
rect 28264 -11266 28266 -11214
rect 28266 -11266 28318 -11214
rect 28318 -11266 28320 -11214
rect 28264 -11268 28320 -11266
rect 33989 -11105 34051 -11101
rect 33989 -11157 34051 -11105
rect 32878 -11291 32950 -11234
rect 33111 -11216 33167 -11212
rect 33111 -11268 33164 -11216
rect 33164 -11268 33167 -11216
rect 27998 -12175 28058 -12117
rect 38833 -11106 38894 -11102
rect 38833 -11158 38894 -11106
rect 37956 -11269 38014 -11213
rect 32888 -12119 32944 -12116
rect 32888 -12171 32889 -12119
rect 32889 -12171 32941 -12119
rect 32941 -12171 32944 -12119
rect 32888 -12173 32944 -12171
rect 42616 -12824 42784 -12656
rect 4893 -13902 4956 -13899
rect 4893 -13955 4956 -13902
rect 3802 -14091 3874 -14035
rect 4035 -14015 4092 -14013
rect 4035 -14067 4037 -14015
rect 4037 -14067 4089 -14015
rect 4089 -14067 4092 -14015
rect 4035 -14070 4092 -14067
rect 3181 -14908 3257 -14903
rect 3181 -14976 3185 -14908
rect 3185 -14976 3254 -14908
rect 3254 -14976 3257 -14908
rect 3181 -14978 3257 -14976
rect 3681 -14983 3746 -14907
rect 9772 -13901 9834 -13898
rect 9772 -13954 9834 -13901
rect 8648 -14091 8720 -14035
rect 8879 -14013 8939 -14011
rect 8879 -14067 8882 -14013
rect 8882 -14067 8937 -14013
rect 8937 -14067 8939 -14013
rect 8879 -14069 8939 -14067
rect 8578 -14919 8636 -14917
rect 8578 -14971 8581 -14919
rect 8581 -14971 8633 -14919
rect 8633 -14971 8636 -14919
rect 8578 -14973 8636 -14971
rect 14580 -13905 14645 -13901
rect 14580 -13957 14645 -13905
rect 13494 -14092 13566 -14035
rect 13725 -14014 13784 -14012
rect 13725 -14067 13727 -14014
rect 13727 -14067 13782 -14014
rect 13782 -14067 13784 -14014
rect 13725 -14069 13784 -14067
rect 13509 -14918 13568 -14916
rect 13509 -14971 13512 -14918
rect 13512 -14971 13567 -14918
rect 13567 -14971 13568 -14918
rect 13509 -14973 13568 -14971
rect 19458 -13906 19521 -13902
rect 19458 -13958 19521 -13906
rect 18340 -14090 18412 -14033
rect 18572 -14013 18630 -14011
rect 18572 -14068 18630 -14013
rect 18252 -14921 18316 -14917
rect 18252 -14974 18256 -14921
rect 18256 -14974 18312 -14921
rect 18312 -14974 18316 -14921
rect 18252 -14979 18316 -14974
rect 24269 -13903 24334 -13899
rect 24269 -13956 24334 -13903
rect 23186 -14092 23258 -14036
rect 23417 -14015 23477 -14013
rect 23417 -14068 23419 -14015
rect 23419 -14068 23474 -14015
rect 23474 -14068 23477 -14015
rect 23417 -14070 23477 -14068
rect 23191 -14913 23254 -14909
rect 23191 -14971 23196 -14913
rect 23196 -14971 23251 -14913
rect 23251 -14971 23254 -14913
rect 23191 -14974 23254 -14971
rect 29145 -13905 29206 -13902
rect 29145 -13958 29206 -13905
rect 28032 -14093 28104 -14037
rect 28263 -14013 28321 -14012
rect 28263 -14067 28264 -14013
rect 28264 -14067 28320 -14013
rect 28320 -14067 28321 -14013
rect 28263 -14068 28321 -14067
rect 33989 -13905 34051 -13901
rect 33989 -13957 34051 -13905
rect 32878 -14093 32950 -14037
rect 33110 -14014 33166 -14012
rect 33110 -14067 33112 -14014
rect 33112 -14067 33164 -14014
rect 33164 -14067 33166 -14014
rect 33110 -14069 33166 -14067
rect 27997 -14972 28062 -14916
rect 38833 -13906 38894 -13902
rect 38833 -13958 38894 -13906
rect 37953 -14068 38013 -14012
rect 32866 -14918 32938 -14916
rect 32866 -14973 32868 -14918
rect 32868 -14973 32936 -14918
rect 32936 -14973 32938 -14918
rect 32866 -14974 32938 -14973
rect 42616 -15624 42784 -15456
rect 4893 -16702 4956 -16699
rect 4893 -16755 4956 -16702
rect 3802 -16891 3874 -16835
rect 4034 -16815 4090 -16812
rect 4034 -16867 4036 -16815
rect 4036 -16867 4088 -16815
rect 4088 -16867 4090 -16815
rect 4034 -16868 4090 -16867
rect 3692 -17783 3760 -17707
rect 9772 -16701 9834 -16698
rect 9772 -16754 9834 -16701
rect 8648 -16892 8720 -16836
rect 8879 -16815 8938 -16812
rect 8879 -16867 8882 -16815
rect 8882 -16867 8934 -16815
rect 8934 -16867 8938 -16815
rect 8879 -16870 8938 -16867
rect 8570 -17720 8630 -17717
rect 8570 -17772 8572 -17720
rect 8572 -17772 8626 -17720
rect 8626 -17772 8630 -17720
rect 8570 -17775 8630 -17772
rect 14580 -16705 14645 -16701
rect 14580 -16757 14645 -16705
rect 13494 -16891 13566 -16835
rect 13726 -16814 13785 -16812
rect 13726 -16867 13728 -16814
rect 13728 -16867 13783 -16814
rect 13783 -16867 13785 -16814
rect 13726 -16869 13785 -16867
rect 19458 -16706 19521 -16702
rect 19458 -16758 19521 -16706
rect 18340 -16892 18412 -16836
rect 18572 -16814 18630 -16810
rect 18572 -16868 18573 -16814
rect 18573 -16868 18627 -16814
rect 18627 -16868 18630 -16814
rect 18572 -16869 18630 -16868
rect 13505 -17717 13561 -17715
rect 13505 -17769 13507 -17717
rect 13507 -17769 13559 -17717
rect 13559 -17769 13561 -17717
rect 13505 -17771 13561 -17769
rect 18250 -17717 18318 -17715
rect 18250 -17773 18253 -17717
rect 18253 -17773 18315 -17717
rect 18315 -17773 18318 -17717
rect 18250 -17776 18318 -17773
rect 24269 -16703 24334 -16699
rect 24269 -16756 24334 -16703
rect 23186 -16893 23258 -16837
rect 23415 -16814 23478 -16811
rect 23415 -16867 23419 -16814
rect 23419 -16867 23475 -16814
rect 23475 -16867 23478 -16814
rect 23415 -16870 23478 -16867
rect 23191 -17714 23251 -17712
rect 23191 -17775 23197 -17714
rect 23197 -17775 23250 -17714
rect 23250 -17775 23251 -17714
rect 23191 -17778 23251 -17775
rect 29145 -16705 29206 -16702
rect 29145 -16758 29206 -16705
rect 28032 -16893 28104 -16837
rect 28265 -16814 28323 -16811
rect 28265 -16866 28267 -16814
rect 28267 -16866 28320 -16814
rect 28320 -16866 28323 -16814
rect 28265 -16867 28323 -16866
rect 27999 -17716 28060 -17712
rect 27999 -17769 28060 -17716
rect 33989 -16705 34051 -16701
rect 33989 -16757 34051 -16705
rect 32878 -16893 32950 -16835
rect 33109 -16815 33167 -16813
rect 33109 -16867 33112 -16815
rect 33112 -16867 33165 -16815
rect 33165 -16867 33167 -16815
rect 33109 -16870 33167 -16867
rect 38833 -16706 38894 -16702
rect 38833 -16758 38894 -16706
rect 37953 -16870 38015 -16808
rect 32868 -17775 32935 -17715
rect 42616 -18424 42784 -18256
rect 4893 -19502 4956 -19499
rect 4893 -19555 4956 -19502
rect 4034 -19615 4091 -19613
rect 4034 -19668 4036 -19615
rect 4036 -19668 4089 -19615
rect 4089 -19668 4091 -19615
rect 4034 -19669 4091 -19668
rect 3696 -20583 3752 -20507
rect 9772 -19501 9834 -19498
rect 9772 -19554 9834 -19501
rect 8881 -19614 8939 -19612
rect 8881 -19666 8882 -19614
rect 8882 -19666 8936 -19614
rect 8936 -19666 8939 -19614
rect 8881 -19668 8939 -19666
rect 8563 -20518 8625 -20514
rect 8563 -20570 8568 -20518
rect 8568 -20570 8620 -20518
rect 8620 -20570 8625 -20518
rect 8563 -20573 8625 -20570
rect 14580 -19505 14645 -19501
rect 14580 -19557 14645 -19505
rect 13727 -19614 13784 -19612
rect 13727 -19666 13729 -19614
rect 13729 -19666 13781 -19614
rect 13781 -19666 13784 -19614
rect 13727 -19668 13784 -19666
rect 19458 -19506 19521 -19502
rect 19458 -19558 19521 -19506
rect 18573 -19669 18630 -19613
rect 13513 -20518 13571 -20515
rect 13513 -20570 13515 -20518
rect 13515 -20570 13568 -20518
rect 13568 -20570 13571 -20518
rect 13513 -20571 13571 -20570
rect 18251 -20521 18315 -20518
rect 18251 -20577 18254 -20521
rect 18254 -20577 18312 -20521
rect 18312 -20577 18315 -20521
rect 18251 -20580 18315 -20577
rect 24269 -19503 24334 -19499
rect 24269 -19556 24334 -19503
rect 23417 -19615 23476 -19612
rect 23417 -19667 23419 -19615
rect 23419 -19667 23474 -19615
rect 23474 -19667 23476 -19615
rect 23417 -19669 23476 -19667
rect 23193 -20517 23253 -20514
rect 23193 -20574 23198 -20517
rect 23198 -20574 23250 -20517
rect 23250 -20574 23253 -20517
rect 23193 -20577 23253 -20574
rect 29145 -19505 29206 -19502
rect 29145 -19558 29206 -19505
rect 28262 -19614 28319 -19612
rect 28262 -19667 28263 -19614
rect 28263 -19667 28318 -19614
rect 28318 -19667 28319 -19614
rect 28262 -19669 28319 -19667
rect 27998 -20574 28059 -20517
rect 33989 -19505 34051 -19501
rect 33989 -19557 34051 -19505
rect 33108 -19614 33170 -19611
rect 33108 -19668 33111 -19614
rect 33111 -19668 33166 -19614
rect 33166 -19668 33170 -19614
rect 33108 -19670 33170 -19668
rect 32869 -20574 32932 -20517
rect 42616 -21224 42785 -21056
<< metal3 >>
rect 3686 2492 3762 2502
rect 3686 2436 3696 2492
rect 3752 2436 3762 2492
rect 3686 2426 3762 2436
rect 8558 2492 8634 2502
rect 8558 2436 8568 2492
rect 8624 2436 8634 2492
rect 8558 2426 8634 2436
rect 13486 2494 13562 2504
rect 13486 2438 13496 2494
rect 13552 2438 13562 2494
rect 13486 2428 13562 2438
rect 18246 2491 18322 2501
rect 18246 2435 18256 2491
rect 18312 2435 18322 2491
rect 18246 2425 18322 2435
rect 23174 2492 23250 2502
rect 23174 2436 23184 2492
rect 23240 2436 23250 2492
rect 23174 2426 23250 2436
rect 27987 2497 28069 2509
rect 27987 2441 28000 2497
rect 28056 2441 28069 2497
rect 27987 2429 28069 2441
rect 32858 2464 32939 2476
rect 32858 2408 32872 2464
rect 32928 2408 32939 2464
rect 32858 2394 32939 2408
rect 23370 1301 23497 1314
rect 13688 1278 13804 1299
rect 13688 1203 13716 1278
rect 13780 1203 13804 1278
rect 13688 1181 13804 1203
rect 18536 1257 18648 1264
rect 18536 1185 18562 1257
rect 18631 1185 18648 1257
rect 23370 1223 23403 1301
rect 23468 1223 23497 1301
rect 23370 1196 23497 1223
rect 28247 1291 28370 1304
rect 28247 1218 28271 1291
rect 28344 1218 28370 1291
rect 28247 1192 28370 1218
rect 33065 1262 33188 1274
rect 33065 1202 33095 1262
rect 33156 1202 33188 1262
rect 18536 1166 18648 1185
rect 33065 1176 33188 1202
rect 6693 888 6807 894
rect 6693 819 6718 888
rect 6790 880 6807 888
rect 6790 876 8945 880
rect 6790 819 8856 876
rect 6693 813 8856 819
rect 8928 813 8945 876
rect 6693 808 8945 813
rect 6693 804 6807 808
rect 3998 537 4115 539
rect 3998 480 4029 537
rect 4093 480 4115 537
rect 3998 448 4115 480
rect 4010 -13 4115 -1
rect 3460 -37 3919 -28
rect 3460 -93 3802 -37
rect 3874 -93 3919 -37
rect 4010 -69 4033 -13
rect 4092 -69 4115 -13
rect 8859 -12 8951 -8
rect 4010 -78 4115 -69
rect 8391 -36 8769 -27
rect 3460 -105 3919 -93
rect 8391 -93 8648 -36
rect 8720 -93 8769 -36
rect 8859 -68 8880 -12
rect 8938 -68 8951 -12
rect 13701 -13 13810 -1
rect 8859 -74 8951 -68
rect 13262 -29 13338 -27
rect 13262 -37 13617 -29
rect 8391 -103 8769 -93
rect 13262 -93 13494 -37
rect 13566 -93 13617 -37
rect 13701 -69 13725 -13
rect 13784 -69 13810 -13
rect 18553 -12 18646 2
rect 13701 -78 13810 -69
rect 18079 -34 18464 -29
rect 3098 -922 3174 -873
rect 3098 -980 3110 -922
rect 3168 -980 3174 -922
rect 3098 -1680 3174 -980
rect 3460 -1680 3536 -105
rect 3672 -907 3794 -884
rect 3672 -983 3696 -907
rect 3774 -983 3794 -907
rect 3672 -1002 3794 -983
rect 8391 -1680 8467 -103
rect 13262 -105 13617 -93
rect 18079 -90 18340 -34
rect 18412 -90 18464 -34
rect 18553 -70 18570 -12
rect 18632 -70 18646 -12
rect 23405 -12 23487 -1
rect 18553 -84 18646 -70
rect 22952 -32 23312 -29
rect 18079 -105 18464 -90
rect 22952 -88 23186 -32
rect 23258 -88 23312 -32
rect 23405 -69 23418 -12
rect 23476 -69 23487 -12
rect 28249 -13 28338 1
rect 23405 -80 23487 -69
rect 27766 -33 28155 -29
rect 22952 -105 23312 -88
rect 27766 -89 28032 -33
rect 28104 -89 28155 -33
rect 28249 -69 28262 -13
rect 28325 -69 28338 -13
rect 33097 -13 33182 -3
rect 28249 -83 28338 -69
rect 32637 -35 32997 -29
rect 27766 -105 28155 -89
rect 32637 -91 32878 -35
rect 32950 -91 32997 -35
rect 33097 -70 33109 -13
rect 33168 -70 33182 -13
rect 33097 -79 33182 -70
rect 37482 -13 38025 -3
rect 37482 -69 37955 -13
rect 38012 -69 38025 -13
rect 37482 -79 38025 -69
rect 32637 -105 32997 -91
rect 8545 -907 8658 -893
rect 8545 -983 8574 -907
rect 8632 -983 8658 -907
rect 8545 -1000 8658 -983
rect 13262 -1680 13338 -105
rect 13469 -916 13581 -896
rect 13469 -974 13505 -916
rect 13567 -974 13581 -916
rect 13469 -998 13581 -974
rect 18079 -1680 18155 -105
rect 18223 -915 18325 -896
rect 18223 -972 18256 -915
rect 18315 -972 18325 -915
rect 18223 -996 18325 -972
rect 22952 -1680 23028 -105
rect 23156 -913 23270 -895
rect 23156 -971 23194 -913
rect 23260 -971 23270 -913
rect 23156 -999 23270 -971
rect 27766 -1680 27842 -105
rect 27975 -915 28081 -898
rect 27975 -975 27999 -915
rect 28058 -975 28081 -915
rect 27975 -1001 28081 -975
rect 32637 -1680 32713 -105
rect 32850 -915 32947 -897
rect 32850 -972 32869 -915
rect 32932 -972 32947 -915
rect 32850 -990 32947 -972
rect 37482 -1680 37558 -79
rect 42560 -1456 42896 1400
rect 42560 -1624 42616 -1456
rect 42784 -1624 42896 -1456
rect 3024 -1848 39032 -1680
rect 4883 -2699 4966 -1848
rect 4883 -2755 4893 -2699
rect 4956 -2755 4966 -2699
rect 4883 -2761 4966 -2755
rect 9762 -2698 9844 -1848
rect 9762 -2754 9772 -2698
rect 9834 -2754 9844 -2698
rect 9762 -2761 9844 -2754
rect 14570 -2701 14655 -1848
rect 14570 -2757 14580 -2701
rect 14645 -2757 14655 -2701
rect 14570 -2761 14655 -2757
rect 19448 -2702 19531 -1848
rect 19448 -2758 19458 -2702
rect 19521 -2758 19531 -2702
rect 19448 -2761 19531 -2758
rect 24259 -2699 24344 -1848
rect 24259 -2756 24269 -2699
rect 24334 -2756 24344 -2699
rect 24259 -2761 24344 -2756
rect 29135 -2702 29216 -1848
rect 29135 -2758 29145 -2702
rect 29206 -2758 29216 -2702
rect 33979 -2701 34061 -1848
rect 33979 -2757 33989 -2701
rect 34051 -2757 34061 -2701
rect 33979 -2761 34061 -2757
rect 38823 -2702 38903 -1848
rect 38823 -2758 38833 -2702
rect 38894 -2758 38904 -2702
rect 38823 -2761 38904 -2758
rect 4009 -2812 4115 -2806
rect 3462 -2835 3924 -2828
rect 3462 -2891 3802 -2835
rect 3874 -2891 3924 -2835
rect 4009 -2868 4035 -2812
rect 4092 -2868 4115 -2812
rect 8860 -2812 8959 -2807
rect 4009 -2875 4115 -2868
rect 8391 -2837 8768 -2828
rect 3462 -2905 3924 -2891
rect 8391 -2893 8648 -2837
rect 8720 -2893 8768 -2837
rect 8860 -2870 8879 -2812
rect 8938 -2870 8959 -2812
rect 13704 -2812 13805 -2804
rect 8860 -2876 8959 -2870
rect 13261 -2835 13615 -2828
rect 8391 -2905 8768 -2893
rect 13261 -2892 13494 -2835
rect 13566 -2892 13615 -2835
rect 13704 -2869 13725 -2812
rect 13784 -2869 13805 -2812
rect 18558 -2812 18642 -2798
rect 13704 -2882 13805 -2869
rect 18080 -2835 18461 -2828
rect 13261 -2905 13615 -2892
rect 18080 -2891 18340 -2835
rect 18412 -2891 18461 -2835
rect 18558 -2870 18570 -2812
rect 18629 -2870 18642 -2812
rect 23402 -2813 23491 -2796
rect 18558 -2878 18642 -2870
rect 22951 -2834 23305 -2828
rect 18080 -2905 18461 -2891
rect 22951 -2890 23186 -2834
rect 23258 -2890 23305 -2834
rect 23402 -2870 23416 -2813
rect 23475 -2870 23491 -2813
rect 28246 -2810 28340 -2801
rect 23402 -2883 23491 -2870
rect 27767 -2834 28150 -2828
rect 22951 -2905 23305 -2890
rect 27767 -2890 28032 -2834
rect 28104 -2890 28150 -2834
rect 28246 -2868 28265 -2810
rect 28322 -2868 28340 -2810
rect 33092 -2813 33180 -2801
rect 28246 -2881 28340 -2868
rect 32639 -2832 33005 -2828
rect 27767 -2905 28150 -2890
rect 32639 -2889 32878 -2832
rect 32950 -2889 33005 -2832
rect 33092 -2869 33110 -2813
rect 33166 -2869 33180 -2813
rect 33092 -2880 33180 -2869
rect 37455 -2834 37847 -2828
rect 32639 -2905 33005 -2889
rect 37455 -2892 37724 -2834
rect 37796 -2892 37847 -2834
rect 37455 -2905 37847 -2892
rect 3082 -3720 3158 -3688
rect 3082 -3780 3092 -3720
rect 3151 -3780 3158 -3720
rect 3082 -4480 3158 -3780
rect 3462 -4480 3538 -2905
rect 3655 -3707 3779 -3692
rect 3655 -3783 3687 -3707
rect 3755 -3783 3779 -3707
rect 3655 -3800 3779 -3783
rect 8391 -4480 8467 -2905
rect 8539 -3707 8643 -3693
rect 8539 -3783 8568 -3707
rect 8628 -3783 8643 -3707
rect 8539 -3797 8643 -3783
rect 13261 -4480 13337 -2905
rect 13472 -3714 13586 -3692
rect 13472 -3774 13507 -3714
rect 13570 -3774 13586 -3714
rect 13472 -3803 13586 -3774
rect 18080 -4480 18156 -2905
rect 18233 -3716 18335 -3695
rect 18233 -3777 18259 -3716
rect 18323 -3777 18335 -3716
rect 18233 -3801 18335 -3777
rect 22951 -4480 23027 -2905
rect 23155 -3718 23270 -3699
rect 23155 -3774 23194 -3718
rect 23253 -3774 23270 -3718
rect 23155 -3796 23270 -3774
rect 27767 -4480 27843 -2905
rect 27965 -3714 28068 -3696
rect 27965 -3772 27990 -3714
rect 28052 -3772 28068 -3714
rect 27965 -3796 28068 -3772
rect 32639 -4480 32715 -2905
rect 32843 -3714 32940 -3695
rect 32843 -3774 32869 -3714
rect 32932 -3774 32940 -3714
rect 32843 -3788 32940 -3774
rect 37455 -4480 37531 -2905
rect 42560 -4256 42896 -1624
rect 42560 -4424 42616 -4256
rect 42784 -4424 42896 -4256
rect 3024 -4648 39032 -4480
rect 4883 -5499 4966 -4648
rect 4883 -5555 4893 -5499
rect 4956 -5555 4966 -5499
rect 4883 -5561 4966 -5555
rect 9762 -5498 9844 -4648
rect 9762 -5554 9772 -5498
rect 9834 -5554 9844 -5498
rect 9762 -5561 9844 -5554
rect 14570 -5501 14655 -4648
rect 14570 -5557 14580 -5501
rect 14645 -5557 14655 -5501
rect 14570 -5561 14655 -5557
rect 19448 -5502 19531 -4648
rect 19448 -5558 19458 -5502
rect 19521 -5558 19531 -5502
rect 19448 -5561 19531 -5558
rect 24259 -5499 24344 -4648
rect 24259 -5556 24269 -5499
rect 24334 -5556 24344 -5499
rect 24259 -5561 24344 -5556
rect 29135 -5502 29216 -4648
rect 29135 -5558 29145 -5502
rect 29206 -5558 29216 -5502
rect 33979 -5501 34061 -4648
rect 33979 -5557 33989 -5501
rect 34051 -5557 34061 -5501
rect 33979 -5561 34061 -5557
rect 38823 -5502 38903 -4648
rect 38823 -5558 38833 -5502
rect 38894 -5558 38904 -5502
rect 38823 -5561 38904 -5558
rect 4015 -5612 4108 -5609
rect 3459 -5637 3917 -5629
rect 3459 -5693 3802 -5637
rect 3874 -5693 3917 -5637
rect 4015 -5668 4035 -5612
rect 4091 -5668 4108 -5612
rect 8860 -5613 8955 -5608
rect 4015 -5675 4108 -5668
rect 8389 -5632 8774 -5627
rect 3459 -5705 3917 -5693
rect 8389 -5690 8648 -5632
rect 8720 -5690 8774 -5632
rect 8860 -5670 8878 -5613
rect 8937 -5670 8955 -5613
rect 13701 -5613 13802 -5602
rect 8860 -5674 8955 -5670
rect 13240 -5635 13620 -5627
rect 8389 -5705 8774 -5690
rect 13240 -5692 13494 -5635
rect 13566 -5692 13620 -5635
rect 13701 -5669 13725 -5613
rect 13783 -5669 13802 -5613
rect 18556 -5607 18645 -5598
rect 13701 -5679 13802 -5669
rect 18078 -5634 18462 -5627
rect 13240 -5705 13620 -5692
rect 18078 -5691 18340 -5634
rect 18412 -5691 18462 -5634
rect 18556 -5671 18569 -5607
rect 18634 -5671 18645 -5607
rect 23404 -5610 23490 -5601
rect 18556 -5682 18645 -5671
rect 22950 -5634 23306 -5627
rect 18078 -5705 18462 -5691
rect 22950 -5691 23186 -5634
rect 23258 -5691 23306 -5634
rect 23404 -5671 23416 -5610
rect 23478 -5671 23490 -5610
rect 28251 -5611 28335 -5601
rect 23404 -5683 23490 -5671
rect 27763 -5634 28155 -5628
rect 22950 -5705 23306 -5691
rect 27763 -5691 28032 -5634
rect 28104 -5691 28155 -5634
rect 28251 -5668 28264 -5611
rect 28323 -5668 28335 -5611
rect 33096 -5611 33179 -5606
rect 28251 -5683 28335 -5668
rect 32639 -5634 33000 -5627
rect 27763 -5705 28155 -5691
rect 32639 -5691 32878 -5634
rect 32950 -5691 33000 -5634
rect 33096 -5669 33109 -5611
rect 33169 -5669 33179 -5611
rect 33096 -5679 33179 -5669
rect 37454 -5612 38029 -5602
rect 37454 -5668 37956 -5612
rect 38014 -5668 38029 -5612
rect 37454 -5678 38029 -5668
rect 32639 -5705 33000 -5691
rect 3077 -6512 3154 -6465
rect 3077 -6569 3087 -6512
rect 3146 -6569 3154 -6512
rect 3077 -7280 3154 -6569
rect 3459 -7280 3535 -5705
rect 3660 -6507 3762 -6493
rect 3660 -6583 3691 -6507
rect 3750 -6583 3762 -6507
rect 3660 -6600 3762 -6583
rect 8389 -7280 8465 -5705
rect 8529 -6507 8634 -6496
rect 8529 -6583 8565 -6507
rect 8624 -6583 8634 -6507
rect 8529 -6597 8634 -6583
rect 13240 -7280 13316 -5705
rect 13470 -6513 13579 -6495
rect 13470 -6573 13506 -6513
rect 13569 -6573 13579 -6513
rect 13470 -6597 13579 -6573
rect 18079 -7280 18155 -5705
rect 18230 -6517 18333 -6492
rect 18230 -6577 18253 -6517
rect 18318 -6577 18333 -6517
rect 18230 -6599 18333 -6577
rect 22950 -7280 23026 -5705
rect 23153 -6516 23268 -6495
rect 23153 -6572 23194 -6516
rect 23252 -6572 23268 -6516
rect 23153 -6597 23268 -6572
rect 27763 -7280 27839 -5705
rect 27963 -6515 28073 -6494
rect 27963 -6576 27985 -6515
rect 28045 -6576 28073 -6515
rect 27963 -6597 28073 -6576
rect 32639 -7280 32715 -5705
rect 32851 -6517 32944 -6500
rect 32851 -6573 32870 -6517
rect 32933 -6573 32944 -6517
rect 32851 -6588 32944 -6573
rect 37454 -7280 37530 -5678
rect 42560 -7056 42896 -4424
rect 42560 -7224 42616 -7056
rect 42784 -7224 42896 -7056
rect 3024 -7448 39032 -7280
rect 3459 -7449 3535 -7448
rect 4883 -8299 4966 -7448
rect 4883 -8355 4893 -8299
rect 4956 -8355 4966 -8299
rect 4883 -8361 4966 -8355
rect 9762 -7498 9845 -7448
rect 9762 -8298 9844 -7498
rect 9762 -8354 9772 -8298
rect 9834 -8354 9844 -8298
rect 9762 -8361 9844 -8354
rect 14570 -8301 14655 -7448
rect 14570 -8357 14580 -8301
rect 14645 -8357 14655 -8301
rect 14570 -8361 14655 -8357
rect 19448 -7488 19533 -7448
rect 19448 -8302 19531 -7488
rect 19448 -8358 19458 -8302
rect 19521 -8358 19531 -8302
rect 19448 -8361 19531 -8358
rect 24259 -8299 24344 -7448
rect 27763 -7449 27839 -7448
rect 24259 -8356 24269 -8299
rect 24334 -8356 24344 -8299
rect 24259 -8361 24344 -8356
rect 29135 -7483 29220 -7448
rect 33979 -7481 34064 -7448
rect 29135 -8302 29216 -7483
rect 29135 -8358 29145 -8302
rect 29206 -8358 29216 -8302
rect 33979 -8301 34061 -7481
rect 33979 -8357 33989 -8301
rect 34051 -8357 34061 -8301
rect 33979 -8361 34061 -8357
rect 38823 -7483 38908 -7448
rect 38823 -8302 38903 -7483
rect 38823 -8358 38833 -8302
rect 38894 -8358 38904 -8302
rect 38823 -8361 38904 -8358
rect 4013 -8413 4113 -8406
rect 3463 -8434 3920 -8429
rect 3463 -8493 3802 -8434
rect 3874 -8493 3920 -8434
rect 4013 -8469 4034 -8413
rect 4091 -8469 4113 -8413
rect 8854 -8411 8968 -8405
rect 4013 -8478 4113 -8469
rect 8391 -8435 8774 -8427
rect 3463 -8505 3920 -8493
rect 8391 -8492 8648 -8435
rect 8720 -8492 8774 -8435
rect 8854 -8471 8878 -8411
rect 8942 -8471 8968 -8411
rect 13705 -8413 13804 -8401
rect 8854 -8481 8968 -8471
rect 13236 -8433 13616 -8427
rect 8391 -8505 8774 -8492
rect 13236 -8491 13494 -8433
rect 13566 -8491 13616 -8433
rect 13705 -8469 13726 -8413
rect 13782 -8469 13804 -8413
rect 18550 -8412 18647 -8398
rect 13705 -8478 13804 -8469
rect 18078 -8433 18464 -8427
rect 13236 -8505 13616 -8491
rect 18078 -8491 18340 -8433
rect 18412 -8491 18464 -8433
rect 18078 -8505 18464 -8491
rect 18550 -8470 18571 -8412
rect 18629 -8470 18647 -8412
rect 23405 -8406 23490 -8393
rect 18550 -8493 18647 -8470
rect 22951 -8434 23310 -8427
rect 22951 -8491 23186 -8434
rect 23258 -8491 23310 -8434
rect 23405 -8471 23416 -8406
rect 23479 -8471 23490 -8406
rect 28247 -8411 28343 -8401
rect 23405 -8481 23490 -8471
rect 27768 -8433 28156 -8427
rect 22951 -8505 23310 -8491
rect 27768 -8492 28032 -8433
rect 28104 -8492 28156 -8433
rect 28247 -8469 28262 -8411
rect 28323 -8469 28343 -8411
rect 33093 -8413 33183 -8403
rect 28247 -8487 28343 -8469
rect 32636 -8434 33000 -8427
rect 27768 -8505 28156 -8492
rect 32636 -8490 32878 -8434
rect 32950 -8490 33000 -8434
rect 33093 -8471 33107 -8413
rect 33166 -8471 33183 -8413
rect 33093 -8484 33183 -8471
rect 37455 -8413 38023 -8403
rect 37455 -8469 37955 -8413
rect 38013 -8469 38023 -8413
rect 37455 -8479 38023 -8469
rect 32636 -8505 33000 -8490
rect 3291 -9400 3367 -9390
rect 3291 -9464 3298 -9400
rect 3362 -9464 3367 -9400
rect 3291 -10080 3367 -9464
rect 3463 -10080 3539 -8505
rect 3670 -9317 3776 -9299
rect 3670 -9373 3696 -9317
rect 3752 -9373 3776 -9317
rect 3670 -9397 3776 -9373
rect 8391 -10080 8467 -8505
rect 8529 -9307 8645 -9296
rect 8529 -9383 8566 -9307
rect 8627 -9383 8645 -9307
rect 8529 -9402 8645 -9383
rect 13236 -10080 13312 -8505
rect 13467 -9314 13579 -9296
rect 13467 -9373 13505 -9314
rect 13570 -9373 13579 -9314
rect 13467 -9399 13579 -9373
rect 18078 -10080 18154 -8505
rect 18226 -9317 18333 -9296
rect 18226 -9376 18252 -9317
rect 18318 -9376 18333 -9317
rect 18226 -9396 18333 -9376
rect 22951 -10080 23027 -8505
rect 23153 -9314 23265 -9295
rect 23153 -9373 23194 -9314
rect 23252 -9373 23265 -9314
rect 23153 -9397 23265 -9373
rect 27768 -10080 27844 -8505
rect 27968 -9317 28077 -9293
rect 27968 -9375 27993 -9317
rect 28053 -9375 28077 -9317
rect 27968 -9397 28077 -9375
rect 32636 -10080 32712 -8505
rect 32853 -9316 32946 -9300
rect 32853 -9374 32867 -9316
rect 32933 -9374 32946 -9316
rect 32853 -9387 32946 -9374
rect 37455 -10080 37531 -8479
rect 42560 -9856 42896 -7224
rect 42560 -10024 42616 -9856
rect 42784 -10024 42896 -9856
rect 3192 -10248 39032 -10080
rect 3463 -10249 3539 -10248
rect 4883 -11099 4966 -10248
rect 4883 -11155 4893 -11099
rect 4956 -11155 4966 -11099
rect 4883 -11161 4966 -11155
rect 9762 -10298 9845 -10248
rect 9762 -11098 9844 -10298
rect 9762 -11154 9772 -11098
rect 9834 -11154 9844 -11098
rect 9762 -11161 9844 -11154
rect 14570 -11101 14655 -10248
rect 14570 -11157 14580 -11101
rect 14645 -11157 14655 -11101
rect 14570 -11161 14655 -11157
rect 19448 -10288 19533 -10248
rect 19448 -11102 19531 -10288
rect 19448 -11158 19458 -11102
rect 19521 -11158 19531 -11102
rect 19448 -11161 19531 -11158
rect 24259 -11099 24344 -10248
rect 24259 -11156 24269 -11099
rect 24334 -11156 24344 -11099
rect 24259 -11161 24344 -11156
rect 29135 -10283 29220 -10248
rect 33979 -10281 34064 -10248
rect 29135 -11102 29216 -10283
rect 29135 -11158 29145 -11102
rect 29206 -11158 29216 -11102
rect 33979 -11101 34061 -10281
rect 33979 -11157 33989 -11101
rect 34051 -11157 34061 -11101
rect 33979 -11161 34061 -11157
rect 38823 -11102 38903 -10248
rect 38823 -11158 38833 -11102
rect 38894 -11158 38904 -11102
rect 38823 -11161 38904 -11158
rect 4013 -11212 4108 -11207
rect 3460 -11232 3924 -11227
rect 3460 -11291 3802 -11232
rect 3874 -11291 3924 -11232
rect 4013 -11268 4035 -11212
rect 4091 -11268 4108 -11212
rect 8855 -11212 8956 -11201
rect 4013 -11277 4108 -11268
rect 8391 -11235 8771 -11227
rect 3460 -11305 3924 -11291
rect 8391 -11291 8648 -11235
rect 8720 -11291 8771 -11235
rect 8855 -11272 8874 -11212
rect 8938 -11272 8956 -11212
rect 13707 -11212 13797 -11202
rect 8855 -11284 8956 -11272
rect 13240 -11233 13617 -11227
rect 8391 -11305 8771 -11291
rect 13240 -11293 13494 -11233
rect 13566 -11293 13617 -11233
rect 13707 -11269 13726 -11212
rect 13782 -11269 13797 -11212
rect 18556 -11210 18647 -11195
rect 13707 -11284 13797 -11269
rect 18082 -11231 18462 -11225
rect 13240 -11305 13617 -11293
rect 18082 -11291 18340 -11231
rect 18412 -11291 18462 -11231
rect 18556 -11270 18571 -11210
rect 18630 -11270 18647 -11210
rect 23405 -11210 23490 -11197
rect 18556 -11284 18647 -11270
rect 22922 -11235 23307 -11226
rect 18082 -11305 18462 -11291
rect 22922 -11293 23186 -11235
rect 23258 -11293 23307 -11235
rect 23405 -11270 23417 -11210
rect 23480 -11270 23490 -11210
rect 28248 -11212 28335 -11204
rect 23405 -11283 23490 -11270
rect 27766 -11234 28148 -11226
rect 22922 -11305 23307 -11293
rect 27766 -11291 28032 -11234
rect 28104 -11291 28148 -11234
rect 28248 -11268 28264 -11212
rect 28320 -11268 28335 -11212
rect 33095 -11212 33179 -11203
rect 28248 -11278 28335 -11268
rect 32638 -11234 32996 -11226
rect 27766 -11305 28148 -11291
rect 32638 -11291 32878 -11234
rect 32950 -11291 32996 -11234
rect 33095 -11268 33111 -11212
rect 33167 -11268 33179 -11212
rect 33095 -11279 33179 -11268
rect 37456 -11213 38024 -11203
rect 37456 -11269 37956 -11213
rect 38014 -11269 38024 -11213
rect 37456 -11279 38024 -11269
rect 32638 -11305 32996 -11291
rect 3182 -12155 3276 -12147
rect 3182 -12228 3197 -12155
rect 3267 -12228 3276 -12155
rect 3182 -12438 3276 -12228
rect 3182 -12880 3277 -12438
rect 3460 -12880 3536 -11305
rect 3665 -12107 3777 -12095
rect 3665 -12183 3688 -12107
rect 3758 -12183 3777 -12107
rect 3665 -12198 3777 -12183
rect 8391 -12880 8467 -11305
rect 8523 -12114 8641 -12093
rect 8523 -12174 8559 -12114
rect 8617 -12174 8641 -12114
rect 8523 -12204 8641 -12174
rect 13240 -12880 13316 -11305
rect 13474 -12116 13574 -12096
rect 13474 -12173 13504 -12116
rect 13564 -12173 13574 -12116
rect 13474 -12192 13574 -12173
rect 18082 -12880 18158 -11305
rect 18221 -12118 18325 -12094
rect 18221 -12177 18249 -12118
rect 18313 -12177 18325 -12118
rect 18221 -12198 18325 -12177
rect 22922 -12880 22998 -11305
rect 23150 -12113 23268 -12095
rect 23150 -12176 23190 -12113
rect 23255 -12176 23268 -12113
rect 23150 -12194 23268 -12176
rect 27766 -12880 27842 -11305
rect 27977 -12117 28074 -12100
rect 27977 -12175 27998 -12117
rect 28058 -12175 28074 -12117
rect 27977 -12195 28074 -12175
rect 32638 -12880 32714 -11305
rect 32865 -12116 32956 -12100
rect 32865 -12173 32888 -12116
rect 32944 -12173 32956 -12116
rect 32865 -12190 32956 -12173
rect 37456 -12880 37532 -11279
rect 42560 -12656 42896 -10024
rect 42560 -12824 42616 -12656
rect 42784 -12824 42896 -12656
rect 3136 -13048 39032 -12880
rect 4883 -13899 4966 -13048
rect 4883 -13955 4893 -13899
rect 4956 -13955 4966 -13899
rect 4883 -13961 4966 -13955
rect 9762 -13898 9844 -13048
rect 9762 -13954 9772 -13898
rect 9834 -13954 9844 -13898
rect 9762 -13961 9844 -13954
rect 14570 -13901 14655 -13048
rect 14570 -13957 14580 -13901
rect 14645 -13957 14655 -13901
rect 14570 -13961 14655 -13957
rect 19448 -13902 19531 -13048
rect 19448 -13958 19458 -13902
rect 19521 -13958 19531 -13902
rect 19448 -13961 19531 -13958
rect 24259 -13899 24344 -13048
rect 24259 -13956 24269 -13899
rect 24334 -13956 24344 -13899
rect 24259 -13961 24344 -13956
rect 29135 -13902 29216 -13048
rect 29135 -13958 29145 -13902
rect 29206 -13958 29216 -13902
rect 33979 -13901 34061 -13048
rect 33979 -13957 33989 -13901
rect 34051 -13957 34061 -13901
rect 33979 -13961 34061 -13957
rect 38823 -13902 38903 -13048
rect 38823 -13958 38833 -13902
rect 38894 -13958 38904 -13902
rect 38823 -13961 38904 -13958
rect 4015 -14013 4108 -14001
rect 3461 -14035 3920 -14028
rect 3461 -14091 3802 -14035
rect 3874 -14091 3920 -14035
rect 4015 -14070 4035 -14013
rect 4092 -14070 4108 -14013
rect 8850 -14011 8968 -13998
rect 4015 -14078 4108 -14070
rect 8392 -14035 8768 -14028
rect 3461 -14105 3920 -14091
rect 8392 -14091 8648 -14035
rect 8720 -14091 8768 -14035
rect 8850 -14069 8879 -14011
rect 8939 -14069 8968 -14011
rect 13707 -14012 13799 -14005
rect 8850 -14080 8968 -14069
rect 13238 -14035 13616 -14029
rect 8392 -14105 8768 -14091
rect 13238 -14092 13494 -14035
rect 13566 -14092 13616 -14035
rect 13707 -14069 13725 -14012
rect 13784 -14069 13799 -14012
rect 18551 -14011 18649 -13996
rect 13707 -14079 13799 -14069
rect 18081 -14033 18462 -14028
rect 13238 -14105 13616 -14092
rect 18081 -14090 18340 -14033
rect 18412 -14090 18462 -14033
rect 18551 -14068 18572 -14011
rect 18630 -14068 18649 -14011
rect 23405 -14013 23488 -14001
rect 18551 -14088 18649 -14068
rect 22950 -14029 23026 -14028
rect 22950 -14036 23308 -14029
rect 18081 -14105 18462 -14090
rect 22950 -14092 23186 -14036
rect 23258 -14092 23308 -14036
rect 23405 -14070 23417 -14013
rect 23477 -14070 23488 -14013
rect 28250 -14012 28333 -14003
rect 23405 -14080 23488 -14070
rect 27767 -14029 27843 -14028
rect 27767 -14037 28151 -14029
rect 22950 -14105 23308 -14092
rect 27767 -14093 28032 -14037
rect 28104 -14093 28151 -14037
rect 28250 -14068 28263 -14012
rect 28321 -14068 28333 -14012
rect 33095 -14012 33178 -14005
rect 28250 -14076 28333 -14068
rect 32638 -14029 32714 -14028
rect 32638 -14037 33000 -14029
rect 27767 -14105 28151 -14093
rect 32638 -14093 32878 -14037
rect 32950 -14093 33000 -14037
rect 33095 -14069 33110 -14012
rect 33166 -14069 33178 -14012
rect 33095 -14078 33178 -14069
rect 37454 -14012 38025 -14002
rect 37454 -14068 37953 -14012
rect 38013 -14068 38025 -14012
rect 37454 -14078 38025 -14068
rect 32638 -14105 33000 -14093
rect 3167 -14903 3269 -14893
rect 3167 -14978 3181 -14903
rect 3257 -14978 3269 -14903
rect 3167 -15680 3269 -14978
rect 3461 -15680 3537 -14105
rect 3656 -14907 3771 -14898
rect 3656 -14983 3681 -14907
rect 3746 -14983 3771 -14907
rect 3656 -14995 3771 -14983
rect 8392 -15680 8468 -14105
rect 8539 -14917 8649 -14896
rect 8539 -14973 8578 -14917
rect 8636 -14973 8649 -14917
rect 8539 -14997 8649 -14973
rect 13238 -15680 13314 -14105
rect 13474 -14916 13578 -14897
rect 13474 -14973 13509 -14916
rect 13568 -14973 13578 -14916
rect 13474 -14991 13578 -14973
rect 18081 -15680 18157 -14105
rect 18227 -14917 18340 -14891
rect 18227 -14979 18252 -14917
rect 18316 -14979 18340 -14917
rect 18227 -15005 18340 -14979
rect 22950 -15680 23026 -14105
rect 23147 -14909 23265 -14892
rect 23147 -14974 23191 -14909
rect 23254 -14974 23265 -14909
rect 23147 -14996 23265 -14974
rect 27767 -15680 27843 -14105
rect 27979 -14916 28076 -14899
rect 27979 -14972 27997 -14916
rect 28062 -14972 28076 -14916
rect 27979 -14989 28076 -14972
rect 32638 -15680 32714 -14105
rect 32845 -14916 32949 -14904
rect 32845 -14974 32866 -14916
rect 32938 -14974 32949 -14916
rect 32845 -14989 32949 -14974
rect 37454 -15680 37530 -14078
rect 42560 -15456 42896 -12824
rect 42560 -15624 42616 -15456
rect 42784 -15624 42896 -15456
rect 3080 -15848 39032 -15680
rect 4883 -16699 4966 -15848
rect 4883 -16755 4893 -16699
rect 4956 -16755 4966 -16699
rect 4883 -16761 4966 -16755
rect 9762 -16698 9844 -15848
rect 13238 -15849 13314 -15848
rect 9762 -16754 9772 -16698
rect 9834 -16754 9844 -16698
rect 9762 -16761 9844 -16754
rect 14570 -16701 14655 -15848
rect 14570 -16757 14580 -16701
rect 14645 -16757 14655 -16701
rect 14570 -16761 14655 -16757
rect 19448 -16702 19531 -15848
rect 19448 -16758 19458 -16702
rect 19521 -16758 19531 -16702
rect 19448 -16761 19531 -16758
rect 24259 -16699 24344 -15848
rect 24259 -16756 24269 -16699
rect 24334 -16756 24344 -16699
rect 24259 -16761 24344 -16756
rect 29135 -16702 29216 -15848
rect 29135 -16758 29145 -16702
rect 29206 -16758 29216 -16702
rect 33979 -16701 34061 -15848
rect 33979 -16757 33989 -16701
rect 34051 -16757 34061 -16701
rect 33979 -16761 34061 -16757
rect 38823 -16702 38903 -15848
rect 38823 -16758 38833 -16702
rect 38894 -16758 38904 -16702
rect 38823 -16761 38904 -16758
rect 37456 -16798 37532 -16797
rect 4018 -16812 4107 -16806
rect 3462 -16829 3538 -16828
rect 3462 -16835 3928 -16829
rect 3462 -16891 3802 -16835
rect 3874 -16891 3928 -16835
rect 4018 -16868 4034 -16812
rect 4090 -16868 4107 -16812
rect 8857 -16812 8959 -16805
rect 4018 -16876 4107 -16868
rect 8390 -16836 8772 -16828
rect 3462 -16905 3928 -16891
rect 8390 -16892 8648 -16836
rect 8720 -16892 8772 -16836
rect 8857 -16870 8879 -16812
rect 8938 -16870 8959 -16812
rect 13710 -16812 13795 -16806
rect 8857 -16879 8959 -16870
rect 13252 -16829 13328 -16828
rect 13252 -16835 13616 -16829
rect 8390 -16905 8772 -16892
rect 13252 -16891 13494 -16835
rect 13566 -16891 13616 -16835
rect 13710 -16869 13726 -16812
rect 13785 -16869 13795 -16812
rect 18558 -16810 18643 -16799
rect 13710 -16881 13795 -16869
rect 18080 -16836 18461 -16828
rect 13252 -16905 13616 -16891
rect 18080 -16892 18340 -16836
rect 18412 -16892 18461 -16836
rect 18558 -16869 18572 -16810
rect 18630 -16869 18643 -16810
rect 23406 -16811 23491 -16801
rect 18558 -16884 18643 -16869
rect 22946 -16829 23022 -16828
rect 22946 -16837 23307 -16829
rect 18080 -16905 18461 -16892
rect 22946 -16893 23186 -16837
rect 23258 -16893 23307 -16837
rect 23406 -16870 23415 -16811
rect 23478 -16870 23491 -16811
rect 28249 -16811 28334 -16804
rect 23406 -16880 23491 -16870
rect 27769 -16829 27845 -16828
rect 27769 -16837 28153 -16829
rect 22946 -16905 23307 -16893
rect 27769 -16893 28032 -16837
rect 28104 -16893 28153 -16837
rect 28249 -16867 28265 -16811
rect 28323 -16867 28334 -16811
rect 33096 -16813 33184 -16801
rect 28249 -16875 28334 -16867
rect 32636 -16829 32712 -16828
rect 32636 -16835 32999 -16829
rect 27769 -16905 28153 -16893
rect 32636 -16893 32878 -16835
rect 32950 -16893 32999 -16835
rect 33096 -16870 33109 -16813
rect 33167 -16870 33184 -16813
rect 33096 -16878 33184 -16870
rect 37456 -16808 38025 -16798
rect 37456 -16870 37953 -16808
rect 38015 -16870 38025 -16808
rect 32636 -16905 32999 -16893
rect 37456 -16880 38025 -16870
rect 3462 -18480 3538 -16905
rect 3664 -17707 3776 -17696
rect 3664 -17783 3692 -17707
rect 3760 -17783 3776 -17707
rect 3664 -17796 3776 -17783
rect 8390 -18480 8466 -16905
rect 8538 -17717 8646 -17693
rect 8538 -17775 8570 -17717
rect 8630 -17775 8646 -17717
rect 8538 -17798 8646 -17775
rect 13252 -18480 13328 -16905
rect 13483 -17715 13572 -17699
rect 13483 -17771 13505 -17715
rect 13561 -17771 13572 -17715
rect 13483 -17793 13572 -17771
rect 18080 -18480 18156 -16905
rect 18221 -17715 18335 -17695
rect 18221 -17776 18250 -17715
rect 18318 -17776 18335 -17715
rect 18221 -17796 18335 -17776
rect 22946 -18480 23022 -16905
rect 23153 -17712 23267 -17694
rect 23153 -17778 23191 -17712
rect 23251 -17778 23267 -17712
rect 23153 -17798 23267 -17778
rect 27769 -18480 27845 -16905
rect 27983 -17712 28077 -17698
rect 27983 -17769 27999 -17712
rect 28060 -17769 28077 -17712
rect 27983 -17787 28077 -17769
rect 32636 -18480 32712 -16905
rect 32850 -17715 32945 -17702
rect 32850 -17775 32868 -17715
rect 32935 -17775 32945 -17715
rect 32850 -17791 32945 -17775
rect 37456 -18480 37532 -16880
rect 42560 -18256 42896 -15624
rect 42560 -18424 42616 -18256
rect 42784 -18424 42896 -18256
rect 3416 -18648 39032 -18480
rect 4883 -19499 4966 -18648
rect 4883 -19555 4893 -19499
rect 4956 -19555 4966 -19499
rect 4883 -19561 4966 -19555
rect 9762 -19498 9844 -18648
rect 9762 -19554 9772 -19498
rect 9834 -19554 9844 -19498
rect 9762 -19561 9844 -19554
rect 14570 -19501 14655 -18648
rect 14570 -19557 14580 -19501
rect 14645 -19557 14655 -19501
rect 14570 -19561 14655 -19557
rect 19448 -19502 19531 -18648
rect 19448 -19558 19458 -19502
rect 19521 -19558 19531 -19502
rect 19448 -19561 19531 -19558
rect 24259 -19499 24344 -18648
rect 24259 -19556 24269 -19499
rect 24334 -19556 24344 -19499
rect 24259 -19561 24344 -19556
rect 29135 -19502 29216 -18648
rect 29135 -19558 29145 -19502
rect 29206 -19558 29216 -19502
rect 33979 -19501 34061 -18648
rect 37456 -18649 37532 -18648
rect 38823 -18649 38903 -18648
rect 33979 -19557 33989 -19501
rect 34051 -19557 34061 -19501
rect 33979 -19561 34061 -19557
rect 4018 -19613 4107 -19608
rect 4018 -19669 4034 -19613
rect 4091 -19669 4107 -19613
rect 4018 -19678 4107 -19669
rect 8862 -19612 8956 -19603
rect 8862 -19668 8881 -19612
rect 8939 -19668 8956 -19612
rect 8862 -19678 8956 -19668
rect 13713 -19612 13794 -19602
rect 13713 -19668 13727 -19612
rect 13784 -19668 13794 -19612
rect 13713 -19676 13794 -19668
rect 18555 -19613 18649 -19595
rect 18555 -19669 18573 -19613
rect 18630 -19669 18649 -19613
rect 18555 -19683 18649 -19669
rect 23404 -19612 23485 -19605
rect 23404 -19669 23417 -19612
rect 23476 -19669 23485 -19612
rect 23404 -19679 23485 -19669
rect 28246 -19612 28338 -19599
rect 28246 -19669 28262 -19612
rect 28319 -19669 28338 -19612
rect 28246 -19681 28338 -19669
rect 33090 -19611 33189 -19600
rect 33090 -19670 33108 -19611
rect 33170 -19670 33189 -19611
rect 33090 -19685 33189 -19670
rect 3664 -20507 3772 -20496
rect 3664 -20583 3696 -20507
rect 3752 -20583 3772 -20507
rect 3664 -20596 3772 -20583
rect 8532 -20514 8651 -20494
rect 8532 -20573 8563 -20514
rect 8625 -20573 8651 -20514
rect 8532 -20601 8651 -20573
rect 13484 -20515 13581 -20501
rect 13484 -20571 13513 -20515
rect 13571 -20571 13581 -20515
rect 13484 -20589 13581 -20571
rect 18223 -20518 18334 -20497
rect 18223 -20580 18251 -20518
rect 18315 -20580 18334 -20518
rect 18223 -20598 18334 -20580
rect 23162 -20514 23270 -20496
rect 23162 -20577 23193 -20514
rect 23253 -20577 23270 -20514
rect 23162 -20597 23270 -20577
rect 27983 -20517 28072 -20496
rect 27983 -20574 27998 -20517
rect 28059 -20574 28072 -20517
rect 27983 -20587 28072 -20574
rect 32859 -20517 32943 -20503
rect 32859 -20574 32869 -20517
rect 32932 -20574 32943 -20517
rect 32859 -20586 32943 -20574
rect 42560 -21056 42896 -18424
rect 42560 -21224 42616 -21056
rect 42785 -21224 42896 -21056
rect 42560 -21392 42896 -21224
<< via3 >>
rect 3696 2436 3752 2492
rect 8568 2436 8624 2492
rect 13496 2438 13552 2494
rect 18256 2435 18312 2491
rect 23184 2436 23240 2492
rect 28000 2441 28056 2497
rect 32872 2408 32928 2464
rect 13716 1203 13780 1278
rect 18562 1185 18631 1257
rect 23403 1223 23468 1301
rect 28271 1218 28344 1291
rect 33095 1202 33156 1262
rect 8856 813 8928 876
rect 4029 480 4093 537
rect 4033 -69 4092 -13
rect 8880 -68 8938 -12
rect 13725 -69 13784 -13
rect 3696 -983 3774 -907
rect 18570 -70 18632 -12
rect 23418 -69 23476 -12
rect 28262 -69 28325 -13
rect 33109 -70 33168 -13
rect 8574 -983 8632 -907
rect 13505 -974 13567 -916
rect 18256 -972 18315 -915
rect 23194 -971 23260 -913
rect 27999 -975 28058 -915
rect 32869 -972 32932 -915
rect 4035 -2868 4092 -2812
rect 8879 -2870 8938 -2812
rect 13725 -2869 13784 -2812
rect 18570 -2870 18629 -2812
rect 23416 -2870 23475 -2813
rect 28265 -2868 28322 -2810
rect 33110 -2869 33166 -2813
rect 3687 -3783 3755 -3707
rect 8568 -3783 8628 -3707
rect 13507 -3774 13570 -3714
rect 18259 -3777 18323 -3716
rect 23194 -3774 23253 -3718
rect 27990 -3772 28052 -3714
rect 32869 -3774 32932 -3714
rect 4035 -5668 4091 -5612
rect 8878 -5670 8937 -5613
rect 13725 -5669 13783 -5613
rect 18569 -5671 18634 -5607
rect 23416 -5671 23478 -5610
rect 28264 -5668 28323 -5611
rect 33109 -5669 33169 -5611
rect 3691 -6583 3750 -6507
rect 8565 -6583 8624 -6507
rect 13506 -6573 13569 -6513
rect 18253 -6577 18318 -6517
rect 23194 -6572 23252 -6516
rect 27985 -6576 28045 -6515
rect 32870 -6573 32933 -6517
rect 4034 -8469 4091 -8413
rect 8878 -8471 8942 -8411
rect 13726 -8469 13782 -8413
rect 18571 -8470 18629 -8412
rect 23416 -8471 23479 -8406
rect 28262 -8469 28323 -8411
rect 33107 -8471 33166 -8413
rect 3696 -9373 3752 -9317
rect 8566 -9383 8627 -9307
rect 13505 -9373 13570 -9314
rect 18252 -9376 18318 -9317
rect 23194 -9373 23252 -9314
rect 27993 -9375 28053 -9317
rect 32867 -9374 32933 -9316
rect 4035 -11268 4091 -11212
rect 8874 -11272 8938 -11212
rect 13726 -11269 13782 -11212
rect 18571 -11270 18630 -11210
rect 23417 -11270 23480 -11210
rect 28264 -11268 28320 -11212
rect 33111 -11268 33167 -11212
rect 3688 -12183 3758 -12107
rect 8559 -12174 8617 -12114
rect 13504 -12173 13564 -12116
rect 18249 -12177 18313 -12118
rect 23190 -12176 23255 -12113
rect 27998 -12175 28058 -12117
rect 32888 -12173 32944 -12116
rect 4035 -14070 4092 -14013
rect 8879 -14069 8939 -14011
rect 13725 -14069 13784 -14012
rect 18572 -14068 18630 -14011
rect 23417 -14070 23477 -14013
rect 28263 -14068 28321 -14012
rect 33110 -14069 33166 -14012
rect 3681 -14983 3746 -14907
rect 8578 -14973 8636 -14917
rect 13509 -14973 13568 -14916
rect 18252 -14979 18316 -14917
rect 23191 -14974 23254 -14909
rect 27997 -14972 28062 -14916
rect 32866 -14974 32938 -14916
rect 4034 -16868 4090 -16812
rect 8879 -16870 8938 -16812
rect 13726 -16869 13785 -16812
rect 18572 -16869 18630 -16810
rect 23415 -16870 23478 -16811
rect 28265 -16867 28323 -16811
rect 33109 -16870 33167 -16813
rect 3692 -17783 3760 -17707
rect 8570 -17775 8630 -17717
rect 13505 -17771 13561 -17715
rect 18250 -17776 18318 -17715
rect 23191 -17778 23251 -17712
rect 27999 -17769 28060 -17712
rect 32868 -17775 32935 -17715
rect 4034 -19669 4091 -19613
rect 8881 -19668 8939 -19612
rect 13727 -19668 13784 -19612
rect 18573 -19669 18630 -19613
rect 23417 -19669 23476 -19612
rect 28262 -19669 28319 -19612
rect 33108 -19670 33170 -19611
rect 3696 -20583 3752 -20507
rect 8563 -20573 8625 -20514
rect 13513 -20571 13571 -20515
rect 18251 -20580 18315 -20518
rect 23193 -20577 23253 -20514
rect 27998 -20574 28059 -20517
rect 32869 -20574 32932 -20517
<< metal4 >>
rect 3640 2492 3808 2632
rect 3640 2436 3696 2492
rect 3752 2436 3808 2492
rect 3640 -907 3808 2436
rect 8512 2492 8680 2632
rect 8512 2436 8568 2492
rect 8624 2436 8680 2492
rect 3640 -983 3696 -907
rect 3774 -983 3808 -907
rect 3640 -3707 3808 -983
rect 3640 -3783 3687 -3707
rect 3755 -3783 3808 -3707
rect 3640 -6507 3808 -3783
rect 3640 -6583 3691 -6507
rect 3750 -6583 3808 -6507
rect 3640 -9317 3808 -6583
rect 3640 -9373 3696 -9317
rect 3752 -9373 3808 -9317
rect 3640 -12107 3808 -9373
rect 3640 -12183 3688 -12107
rect 3758 -12183 3808 -12107
rect 3640 -14907 3808 -12183
rect 3640 -14983 3681 -14907
rect 3746 -14983 3808 -14907
rect 3640 -17707 3808 -14983
rect 3640 -17783 3692 -17707
rect 3760 -17783 3808 -17707
rect 3640 -20507 3808 -17783
rect 3640 -20583 3696 -20507
rect 3752 -20583 3808 -20507
rect 3640 -21224 3808 -20583
rect 3976 537 4144 560
rect 3976 480 4029 537
rect 4093 480 4144 537
rect 3976 -13 4144 480
rect 3976 -69 4033 -13
rect 4092 -69 4144 -13
rect 3976 -2812 4144 -69
rect 3976 -2868 4035 -2812
rect 4092 -2868 4144 -2812
rect 3976 -5612 4144 -2868
rect 3976 -5668 4035 -5612
rect 4091 -5668 4144 -5612
rect 3976 -8413 4144 -5668
rect 3976 -8469 4034 -8413
rect 4091 -8469 4144 -8413
rect 3976 -11212 4144 -8469
rect 3976 -11268 4035 -11212
rect 4091 -11268 4144 -11212
rect 3976 -14013 4144 -11268
rect 3976 -14070 4035 -14013
rect 4092 -14070 4144 -14013
rect 3976 -16812 4144 -14070
rect 3976 -16868 4034 -16812
rect 4090 -16868 4144 -16812
rect 3976 -19613 4144 -16868
rect 3976 -19669 4034 -19613
rect 4091 -19669 4144 -19613
rect 3976 -21224 4144 -19669
rect 8512 -907 8680 2436
rect 13440 2494 13608 2632
rect 13440 2438 13496 2494
rect 13552 2438 13608 2494
rect 8512 -983 8574 -907
rect 8632 -983 8680 -907
rect 8512 -3707 8680 -983
rect 8512 -3783 8568 -3707
rect 8628 -3783 8680 -3707
rect 8512 -6507 8680 -3783
rect 8512 -6583 8565 -6507
rect 8624 -6583 8680 -6507
rect 8512 -9307 8680 -6583
rect 8512 -9383 8566 -9307
rect 8627 -9383 8680 -9307
rect 8512 -12114 8680 -9383
rect 8512 -12174 8559 -12114
rect 8617 -12174 8680 -12114
rect 8512 -14917 8680 -12174
rect 8512 -14973 8578 -14917
rect 8636 -14973 8680 -14917
rect 8512 -17717 8680 -14973
rect 8512 -17775 8570 -17717
rect 8630 -17775 8680 -17717
rect 8512 -20514 8680 -17775
rect 8512 -20573 8563 -20514
rect 8625 -20573 8680 -20514
rect 8512 -21392 8680 -20573
rect 8818 876 8996 1039
rect 8818 813 8856 876
rect 8928 813 8996 876
rect 8818 -12 8996 813
rect 8818 -68 8880 -12
rect 8938 -68 8996 -12
rect 8818 -2812 8996 -68
rect 8818 -2870 8879 -2812
rect 8938 -2870 8996 -2812
rect 8818 -5613 8996 -2870
rect 8818 -5670 8878 -5613
rect 8937 -5670 8996 -5613
rect 8818 -8411 8996 -5670
rect 8818 -8471 8878 -8411
rect 8942 -8471 8996 -8411
rect 8818 -11212 8996 -8471
rect 8818 -11272 8874 -11212
rect 8938 -11272 8996 -11212
rect 8818 -14011 8996 -11272
rect 8818 -14069 8879 -14011
rect 8939 -14069 8996 -14011
rect 8818 -16812 8996 -14069
rect 8818 -16870 8879 -16812
rect 8938 -16870 8996 -16812
rect 8818 -19612 8996 -16870
rect 8818 -19668 8881 -19612
rect 8939 -19668 8996 -19612
rect 8818 -21392 8996 -19668
rect 13440 -916 13608 2438
rect 18200 2491 18368 2632
rect 18200 2435 18256 2491
rect 18312 2435 18368 2491
rect 13440 -974 13505 -916
rect 13567 -974 13608 -916
rect 13440 -3714 13608 -974
rect 13440 -3774 13507 -3714
rect 13570 -3774 13608 -3714
rect 13440 -6513 13608 -3774
rect 13440 -6573 13506 -6513
rect 13569 -6573 13608 -6513
rect 13440 -9314 13608 -6573
rect 13440 -9373 13505 -9314
rect 13570 -9373 13608 -9314
rect 13440 -12116 13608 -9373
rect 13440 -12173 13504 -12116
rect 13564 -12173 13608 -12116
rect 13440 -14916 13608 -12173
rect 13440 -14973 13509 -14916
rect 13568 -14973 13608 -14916
rect 13440 -17715 13608 -14973
rect 13440 -17771 13505 -17715
rect 13561 -17771 13608 -17715
rect 13440 -20515 13608 -17771
rect 13440 -20571 13513 -20515
rect 13571 -20571 13608 -20515
rect 13440 -21336 13608 -20571
rect 13664 1278 13832 1344
rect 13664 1203 13716 1278
rect 13780 1203 13832 1278
rect 13664 952 13832 1203
rect 13664 -13 13833 952
rect 13664 -69 13725 -13
rect 13784 -69 13833 -13
rect 13664 -2812 13833 -69
rect 13664 -2869 13725 -2812
rect 13784 -2869 13833 -2812
rect 13664 -5613 13833 -2869
rect 13664 -5669 13725 -5613
rect 13783 -5669 13833 -5613
rect 13664 -8413 13833 -5669
rect 13664 -8469 13726 -8413
rect 13782 -8469 13833 -8413
rect 13664 -11212 13833 -8469
rect 13664 -11269 13726 -11212
rect 13782 -11269 13833 -11212
rect 13664 -14012 13833 -11269
rect 13664 -14069 13725 -14012
rect 13784 -14069 13833 -14012
rect 13664 -16812 13833 -14069
rect 13664 -16869 13726 -16812
rect 13785 -16869 13833 -16812
rect 13664 -19612 13833 -16869
rect 13664 -19668 13727 -19612
rect 13784 -19668 13833 -19612
rect 13664 -21336 13833 -19668
rect 18200 -915 18368 2435
rect 23128 2492 23296 2632
rect 23128 2436 23184 2492
rect 23240 2436 23296 2492
rect 18200 -972 18256 -915
rect 18315 -972 18368 -915
rect 18200 -3716 18368 -972
rect 18200 -3777 18259 -3716
rect 18323 -3777 18368 -3716
rect 18200 -6517 18368 -3777
rect 18200 -6577 18253 -6517
rect 18318 -6577 18368 -6517
rect 18200 -9317 18368 -6577
rect 18200 -9376 18252 -9317
rect 18318 -9376 18368 -9317
rect 18200 -12118 18368 -9376
rect 18200 -12177 18249 -12118
rect 18313 -12177 18368 -12118
rect 18200 -14917 18368 -12177
rect 18200 -14979 18252 -14917
rect 18316 -14979 18368 -14917
rect 18200 -17715 18368 -14979
rect 18200 -17776 18250 -17715
rect 18318 -17776 18368 -17715
rect 18200 -20518 18368 -17776
rect 18200 -20580 18251 -20518
rect 18315 -20580 18368 -20518
rect 18200 -21336 18368 -20580
rect 18505 1257 18674 1278
rect 18505 1185 18562 1257
rect 18631 1185 18674 1257
rect 18505 -12 18674 1185
rect 18505 -70 18570 -12
rect 18632 -70 18674 -12
rect 18505 -2812 18674 -70
rect 18505 -2870 18570 -2812
rect 18629 -2870 18674 -2812
rect 18505 -5607 18674 -2870
rect 18505 -5671 18569 -5607
rect 18634 -5671 18674 -5607
rect 18505 -8412 18674 -5671
rect 18505 -8470 18571 -8412
rect 18629 -8470 18674 -8412
rect 18505 -11210 18674 -8470
rect 18505 -11270 18571 -11210
rect 18630 -11270 18674 -11210
rect 18505 -14011 18674 -11270
rect 18505 -14068 18572 -14011
rect 18630 -14068 18674 -14011
rect 18505 -16810 18674 -14068
rect 18505 -16869 18572 -16810
rect 18630 -16869 18674 -16810
rect 18505 -19613 18674 -16869
rect 18505 -19669 18573 -19613
rect 18630 -19669 18674 -19613
rect 18505 -21336 18674 -19669
rect 23128 -913 23296 2436
rect 27944 2497 28112 2632
rect 27944 2441 28000 2497
rect 28056 2441 28112 2497
rect 23128 -971 23194 -913
rect 23260 -971 23296 -913
rect 23128 -3718 23296 -971
rect 23128 -3774 23194 -3718
rect 23253 -3774 23296 -3718
rect 23128 -6516 23296 -3774
rect 23128 -6572 23194 -6516
rect 23252 -6572 23296 -6516
rect 23128 -9314 23296 -6572
rect 23128 -9373 23194 -9314
rect 23252 -9373 23296 -9314
rect 23128 -12113 23296 -9373
rect 23128 -12176 23190 -12113
rect 23255 -12176 23296 -12113
rect 23128 -14909 23296 -12176
rect 23128 -14974 23191 -14909
rect 23254 -14974 23296 -14909
rect 23128 -17712 23296 -14974
rect 23128 -17778 23191 -17712
rect 23251 -17778 23296 -17712
rect 23128 -20514 23296 -17778
rect 23128 -20577 23193 -20514
rect 23253 -20577 23296 -20514
rect 23128 -21336 23296 -20577
rect 23352 1301 23520 1344
rect 23352 1223 23403 1301
rect 23468 1223 23520 1301
rect 23352 -12 23520 1223
rect 23352 -69 23418 -12
rect 23476 -69 23520 -12
rect 23352 -2813 23520 -69
rect 23352 -2870 23416 -2813
rect 23475 -2870 23520 -2813
rect 23352 -5610 23520 -2870
rect 23352 -5671 23416 -5610
rect 23478 -5671 23520 -5610
rect 23352 -8406 23520 -5671
rect 23352 -8471 23416 -8406
rect 23479 -8471 23520 -8406
rect 23352 -11210 23520 -8471
rect 23352 -11270 23417 -11210
rect 23480 -11270 23520 -11210
rect 23352 -14013 23520 -11270
rect 23352 -14070 23417 -14013
rect 23477 -14070 23520 -14013
rect 23352 -16811 23520 -14070
rect 23352 -16870 23415 -16811
rect 23478 -16870 23520 -16811
rect 23352 -19612 23520 -16870
rect 23352 -19669 23417 -19612
rect 23476 -19669 23520 -19612
rect 23352 -21336 23520 -19669
rect 27944 -915 28112 2441
rect 32816 2464 32984 2632
rect 32816 2408 32872 2464
rect 32928 2408 32984 2464
rect 27944 -975 27999 -915
rect 28058 -975 28112 -915
rect 27944 -3714 28112 -975
rect 27944 -3772 27990 -3714
rect 28052 -3772 28112 -3714
rect 27944 -6515 28112 -3772
rect 27944 -6576 27985 -6515
rect 28045 -6576 28112 -6515
rect 27944 -9317 28112 -6576
rect 27944 -9375 27993 -9317
rect 28053 -9375 28112 -9317
rect 27944 -12117 28112 -9375
rect 27944 -12175 27998 -12117
rect 28058 -12175 28112 -12117
rect 27944 -14916 28112 -12175
rect 27944 -14972 27997 -14916
rect 28062 -14972 28112 -14916
rect 27944 -17712 28112 -14972
rect 27944 -17769 27999 -17712
rect 28060 -17769 28112 -17712
rect 27944 -20517 28112 -17769
rect 27944 -20574 27998 -20517
rect 28059 -20574 28112 -20517
rect 27944 -21336 28112 -20574
rect 28224 1291 28392 1336
rect 28224 1218 28271 1291
rect 28344 1218 28392 1291
rect 28224 -13 28392 1218
rect 28224 -69 28262 -13
rect 28325 -69 28392 -13
rect 28224 -2810 28392 -69
rect 28224 -2868 28265 -2810
rect 28322 -2868 28392 -2810
rect 28224 -5611 28392 -2868
rect 28224 -5668 28264 -5611
rect 28323 -5668 28392 -5611
rect 28224 -8411 28392 -5668
rect 28224 -8469 28262 -8411
rect 28323 -8469 28392 -8411
rect 28224 -11212 28392 -8469
rect 28224 -11268 28264 -11212
rect 28320 -11268 28392 -11212
rect 28224 -14012 28392 -11268
rect 28224 -14068 28263 -14012
rect 28321 -14068 28392 -14012
rect 28224 -16811 28392 -14068
rect 28224 -16867 28265 -16811
rect 28323 -16867 28392 -16811
rect 28224 -19612 28392 -16867
rect 28224 -19669 28262 -19612
rect 28319 -19669 28392 -19612
rect 28224 -21336 28392 -19669
rect 32816 -915 32984 2408
rect 32816 -972 32869 -915
rect 32932 -972 32984 -915
rect 32816 -3714 32984 -972
rect 32816 -3774 32869 -3714
rect 32932 -3774 32984 -3714
rect 32816 -6517 32984 -3774
rect 32816 -6573 32870 -6517
rect 32933 -6573 32984 -6517
rect 32816 -9316 32984 -6573
rect 32816 -9374 32867 -9316
rect 32933 -9374 32984 -9316
rect 32816 -12116 32984 -9374
rect 32816 -12173 32888 -12116
rect 32944 -12173 32984 -12116
rect 32816 -14916 32984 -12173
rect 32816 -14974 32866 -14916
rect 32938 -14974 32984 -14916
rect 32816 -17715 32984 -14974
rect 32816 -17775 32868 -17715
rect 32935 -17775 32984 -17715
rect 32816 -20517 32984 -17775
rect 32816 -20574 32869 -20517
rect 32932 -20574 32984 -20517
rect 32816 -21392 32984 -20574
rect 33040 1262 33208 1288
rect 33040 1202 33095 1262
rect 33156 1202 33208 1262
rect 33040 -13 33208 1202
rect 33040 -70 33109 -13
rect 33168 -70 33208 -13
rect 33040 -2813 33208 -70
rect 33040 -2869 33110 -2813
rect 33166 -2869 33208 -2813
rect 33040 -5611 33208 -2869
rect 33040 -5669 33109 -5611
rect 33169 -5669 33208 -5611
rect 33040 -8413 33208 -5669
rect 33040 -8471 33107 -8413
rect 33166 -8471 33208 -8413
rect 33040 -11212 33208 -8471
rect 33040 -11268 33111 -11212
rect 33167 -11268 33208 -11212
rect 33040 -14012 33208 -11268
rect 33040 -14069 33110 -14012
rect 33166 -14069 33208 -14012
rect 33040 -16813 33208 -14069
rect 33040 -16870 33109 -16813
rect 33167 -16870 33208 -16813
rect 33040 -19611 33208 -16870
rect 33040 -19670 33108 -19611
rect 33170 -19670 33208 -19611
rect 33040 -21392 33208 -19670
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2506 0 1 -12537
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_1
timestamp 1753044640
transform 1 0 2384 0 -1 -5249
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_2
timestamp 1753044640
transform 1 0 2490 0 1 -18137
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_3
timestamp 1753044640
transform 1 0 2493 0 1 -15337
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_4
timestamp 1753044640
transform 1 0 2490 0 -1 -16449
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_5
timestamp 1753044640
transform 1 0 22038 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_6
timestamp 1753044640
transform 1 0 11286 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_7
timestamp 1753044640
transform 1 0 27078 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_8
timestamp 1753044640
transform 1 0 31726 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_9
timestamp 1753044640
transform 1 0 30606 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2602 0 1 -9737
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_1
timestamp 1753044640
transform 1 0 17278 0 1 1038
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_0 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2403 0 -1 351
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_1
timestamp 1753044640
transform 1 0 2388 0 1 -4137
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_2
timestamp 1753044640
transform 1 0 2403 0 1 -1337
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_3
timestamp 1753044640
transform 1 0 2394 0 -1 -10849
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_4
timestamp 1753044640
transform 1 0 2384 0 1 -6937
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_5
timestamp 1753044640
transform 1 0 2403 0 1 471
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_6
timestamp 1753044640
transform 1 0 2403 0 -1 2159
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_7
timestamp 1753044640
transform 1 0 6022 0 1 471
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_8
timestamp 1753044640
transform 1 0 20918 0 1 1038
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_9
timestamp 1753044640
transform 1 0 12294 0 1 1038
box -86 -86 1206 870
use unit_cell_array  unit_cell_array_0 ~/CS_DAC/Magic_gf180mcuD
timestamp 1754909118
transform 1 0 13288 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_1
timestamp 1754909118
transform 1 0 3596 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_2
timestamp 1754909118
transform 1 0 8442 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_3
timestamp 1754909118
transform 1 0 37518 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_4
timestamp 1754909118
transform 1 0 18134 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_5
timestamp 1754909118
transform 1 0 22980 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_6
timestamp 1754909118
transform 1 0 27826 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_7
timestamp 1754909118
transform 1 0 32672 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_8
timestamp 1754909118
transform 1 0 8442 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_9
timestamp 1754909118
transform 1 0 3596 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_10
timestamp 1754909118
transform 1 0 13288 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_11
timestamp 1754909118
transform 1 0 22980 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_12
timestamp 1754909118
transform 1 0 18134 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_13
timestamp 1754909118
transform 1 0 27826 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_14
timestamp 1754909118
transform 1 0 37518 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_15
timestamp 1754909118
transform 1 0 32672 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_17
timestamp 1754909118
transform 1 0 32672 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_18
timestamp 1754909118
transform 1 0 27826 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_19
timestamp 1754909118
transform 1 0 22980 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_20
timestamp 1754909118
transform 1 0 18134 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_21
timestamp 1754909118
transform 1 0 13288 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_22
timestamp 1754909118
transform 1 0 8442 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_23
timestamp 1754909118
transform 1 0 3596 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_24
timestamp 1754909118
transform 1 0 8442 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_25
timestamp 1754909118
transform 1 0 3596 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_26
timestamp 1754909118
transform 1 0 13288 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_27
timestamp 1754909118
transform 1 0 22980 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_28
timestamp 1754909118
transform 1 0 18134 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_29
timestamp 1754909118
transform 1 0 27826 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_30
timestamp 1754909118
transform 1 0 37518 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_31
timestamp 1754909118
transform 1 0 32672 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_32
timestamp 1754909118
transform 1 0 8442 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_33
timestamp 1754909118
transform 1 0 3596 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_34
timestamp 1754909118
transform 1 0 13288 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_35
timestamp 1754909118
transform 1 0 22980 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_36
timestamp 1754909118
transform 1 0 18134 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_37
timestamp 1754909118
transform 1 0 27826 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_38
timestamp 1754909118
transform 1 0 37518 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_39
timestamp 1754909118
transform 1 0 32672 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_40
timestamp 1754909118
transform 1 0 8442 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_41
timestamp 1754909118
transform 1 0 3596 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_42
timestamp 1754909118
transform 1 0 13288 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_43
timestamp 1754909118
transform 1 0 22980 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_44
timestamp 1754909118
transform 1 0 18134 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_45
timestamp 1754909118
transform 1 0 27826 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_46
timestamp 1754909118
transform 1 0 37518 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_47
timestamp 1754909118
transform 1 0 32672 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_48
timestamp 1754909118
transform 1 0 8442 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_49
timestamp 1754909118
transform 1 0 3596 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_50
timestamp 1754909118
transform 1 0 13288 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_51
timestamp 1754909118
transform 1 0 22980 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_52
timestamp 1754909118
transform 1 0 18134 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_53
timestamp 1754909118
transform 1 0 27826 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_54
timestamp 1754909118
transform 1 0 37518 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_55
timestamp 1754909118
transform 1 0 32672 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_56
timestamp 1754909118
transform 1 0 8442 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_57
timestamp 1754909118
transform 1 0 3596 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_58
timestamp 1754909118
transform 1 0 13288 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_59
timestamp 1754909118
transform 1 0 22980 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_60
timestamp 1754909118
transform 1 0 18134 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_61
timestamp 1754909118
transform 1 0 27826 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_62
timestamp 1754909118
transform 1 0 37518 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_63
timestamp 1754909118
transform 1 0 32672 0 1 -17054
box -12 -1202 4834 691
<< end >>
