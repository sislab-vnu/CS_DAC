magic
tech gf180mcuD
magscale 1 10
timestamp 1756794861
<< metal1 >>
rect 21672 41608 21840 41720
rect 21672 41496 21728 41608
rect 21784 41496 21840 41608
rect -7144 39928 -4624 39929
rect -4256 39928 -4088 39929
rect -9800 39872 -4088 39928
rect -9800 39816 -9744 39872
rect -9688 39816 -4088 39872
rect -9800 39761 -4088 39816
rect -9800 39760 -7127 39761
rect -4872 39760 -4088 39761
rect -4256 18310 -4088 39760
rect -1064 39872 1568 39928
rect -1064 39816 1456 39872
rect 1512 39816 1568 39872
rect -1064 39760 1568 39816
rect -1064 18278 -896 39760
rect 12543 33432 14003 33488
rect 12543 33376 12600 33432
rect 12656 33376 14003 33432
rect 12543 33319 14003 33376
rect 7000 30240 17009 30296
rect 7000 30184 7056 30240
rect 7112 30184 17009 30240
rect 7000 30128 17009 30184
rect 21672 29232 21840 41496
rect 45361 34833 56056 34906
rect 45361 34663 55775 34833
rect 55944 34663 56056 34833
rect 45361 34570 56056 34663
rect 45361 34554 45696 34570
rect 45360 33578 45696 34554
rect 45862 34266 54918 34267
rect 58293 34266 58685 34267
rect 45862 34186 61377 34266
rect 45862 34016 61067 34186
rect 61236 34016 61377 34186
rect 45862 33931 61377 34016
rect 45864 33638 46200 33931
rect 54563 33930 61377 33931
rect 56056 33929 61377 33930
rect 46369 33656 50905 33657
rect 46369 33572 66697 33656
rect 46369 33402 66383 33572
rect 66552 33402 66697 33572
rect 46369 33321 66697 33402
rect 50730 33320 66697 33321
rect 61376 33319 66697 33320
rect 0 29065 39368 29232
rect 0 29064 38914 29065
<< via1 >>
rect 21728 41496 21784 41608
rect -9744 39816 -9688 39872
rect 1456 39816 1512 39872
rect 12600 33376 12656 33432
rect 7056 30184 7112 30240
rect 55775 34663 55944 34833
rect 61067 34016 61236 34186
rect 66383 33402 66552 33572
<< metal2 >>
rect -9800 39872 -9632 41718
rect -9800 39816 -9744 39872
rect -9688 39816 -9632 39872
rect -9800 39760 -9632 39816
rect -3921 39647 -3752 41718
rect 1400 39872 1568 41718
rect 1400 39816 1456 39872
rect 1512 39816 1568 39872
rect 1400 39760 1568 39816
rect -3920 18262 -3752 39647
rect 7000 30240 7168 41718
rect 12543 39983 12711 41718
rect 12543 39704 12712 39983
rect 12543 33432 12711 39704
rect 12543 33376 12600 33432
rect 12656 33376 12711 33432
rect 12543 33319 12711 33376
rect 18088 33095 18256 41718
rect 21672 41608 21840 41720
rect 21672 41496 21728 41608
rect 21784 41496 21840 41608
rect 21672 41384 21840 41496
rect 7000 30184 7056 30240
rect 7112 30184 7168 30240
rect 23632 30352 23800 41718
rect 29232 30856 29400 41718
rect 34832 39732 35000 41718
rect 34831 39207 35000 39732
rect 34832 37605 35000 39207
rect 34831 32200 35000 37605
rect 40432 32872 40600 41718
rect 55664 34833 56056 34906
rect 55664 34663 55775 34833
rect 55944 34663 56056 34833
rect 55664 34570 56056 34663
rect 60928 34186 61377 34266
rect 60928 34016 61067 34186
rect 61236 34016 61377 34186
rect 60928 33929 61377 34016
rect 66248 33572 66697 33656
rect 66248 33402 66383 33572
rect 66552 33402 66697 33572
rect 66248 33319 66697 33402
rect 40480 32865 40561 32872
rect 34831 31976 34999 32200
rect 34831 31808 40558 31976
rect 29232 30688 40486 30856
rect 23632 30184 38864 30352
rect 7000 30128 7168 30184
rect 14440 29904 14478 29913
rect 335 29792 14478 29904
rect 335 29130 503 29792
rect 15344 29680 15401 29928
rect 5935 29568 15401 29680
rect 5935 29057 6103 29568
rect 16240 29456 16298 29910
rect 11535 29344 16298 29456
rect 17192 29344 17249 29969
rect 18032 29456 18089 29931
rect 18984 29909 18985 29929
rect 18928 29680 18985 29909
rect 19824 29792 34103 29904
rect 18928 29568 28503 29680
rect 18032 29344 22902 29456
rect 11535 29187 11703 29344
rect 17135 29120 17304 29344
rect 22735 29133 22902 29344
rect 28335 29157 28503 29568
rect 33935 29134 34103 29792
rect 38696 29736 38864 30184
rect 38696 29568 40560 29736
rect -672 25648 -560 25704
rect -672 25592 -645 25648
rect -589 25592 -560 25648
rect -672 17472 -560 25592
rect -448 22064 -336 22120
rect -448 22008 -422 22064
rect -366 22008 -336 22064
rect -448 16632 -336 22008
rect -674 16576 -336 16632
rect -224 18480 -112 18536
rect -224 18424 -196 18480
rect -140 18424 -112 18480
rect -224 15736 -112 18424
rect -673 15680 -112 15736
rect -224 14896 -110 14923
rect -689 14840 -195 14896
rect -139 14840 -110 14896
rect -224 14809 -110 14840
rect -678 13888 -112 13944
rect -673 12992 -336 13048
rect -672 4144 -560 12125
rect -448 7728 -336 12992
rect -224 11326 -112 13888
rect -224 11270 -202 11326
rect -146 11270 -112 11326
rect -224 11214 -112 11270
rect -448 7672 -416 7728
rect -360 7672 -336 7728
rect -448 7630 -336 7672
rect -672 4088 -644 4144
rect -588 4088 -560 4144
rect -672 4046 -560 4088
<< via2 >>
rect -645 25592 -589 25648
rect 671 25606 727 25662
rect -422 22008 -366 22064
rect 671 22022 727 22078
rect -196 18424 -140 18480
rect 671 18438 727 18494
rect -195 14840 -139 14896
rect 671 14854 727 14910
rect -202 11270 -146 11326
rect 671 11270 727 11326
rect -416 7672 -360 7728
rect 671 7686 727 7742
rect -644 4088 -588 4144
rect 671 4102 727 4158
<< metal3 >>
rect -11033 39634 -6661 39636
rect 49160 39634 55146 39636
rect -11033 37802 55146 39634
rect -11033 37800 51109 37802
rect -11033 37798 -6661 37800
rect -11033 27216 -9199 37798
rect 2139 28952 2363 37800
rect 3248 35401 4089 35504
rect 3248 34775 3327 35401
rect 3994 34775 4089 35401
rect 3248 34663 4089 34775
rect 3539 34408 3764 34663
rect 3539 28948 3763 34408
rect 7739 28056 7963 37800
rect 8791 35402 9632 35504
rect 8791 34776 8907 35402
rect 9574 34776 9632 35402
rect 8791 34663 9632 34776
rect 9139 34507 9364 34663
rect 9139 28000 9363 34507
rect 13339 31361 13563 37800
rect 18939 37755 19163 37800
rect 20750 35402 21591 35503
rect 20750 34776 20850 35402
rect 21517 34776 21591 35402
rect 20750 34662 21591 34776
rect 21075 34379 21300 34662
rect 21075 32368 21299 34379
rect 20705 32148 21299 32368
rect 20705 32144 21018 32148
rect 21075 32092 21299 32148
rect 13339 31136 13971 31361
rect 13339 28056 13563 31136
rect 21074 31087 21299 32092
rect 21074 30616 21298 31087
rect 20339 30392 21298 30616
rect 20339 28916 20563 30392
rect 18939 28280 19163 28397
rect 24539 28280 24763 37800
rect 25674 35404 26515 35505
rect 25674 34778 25772 35404
rect 26439 34778 26515 35404
rect 25674 34664 26515 34778
rect 25939 27999 26163 34664
rect 30139 28280 30363 37800
rect 31248 35399 32089 35505
rect 31248 34773 31321 35399
rect 31988 34773 32089 35399
rect 31248 34664 32089 34773
rect 31539 28248 31763 34664
rect 35739 28280 35963 37800
rect 36848 35400 37689 35505
rect 36848 34774 36928 35400
rect 37595 34774 37689 35400
rect 36848 34664 37689 34774
rect 37139 28275 37363 34664
rect 40655 33666 40881 37800
rect 42055 35392 42897 35504
rect 42055 34776 42168 35392
rect 42785 34776 42897 35392
rect 42055 34664 42897 34776
rect 42280 33682 42504 34664
rect -11033 27124 -4199 27216
rect -11033 26956 -4480 27124
rect -4312 26956 -4199 27124
rect -11033 26880 -4199 26956
rect -11033 20048 -9199 26880
rect 40655 26695 40881 29011
rect 40655 26472 41563 26695
rect 40751 26471 41563 26472
rect -672 25662 784 25718
rect -672 25648 671 25662
rect -672 25592 -645 25648
rect -589 25606 671 25648
rect 727 25606 784 25662
rect -589 25592 784 25606
rect -672 25550 784 25592
rect 41339 25327 41563 26471
rect 42280 26472 42504 29009
rect 53312 27216 55146 37802
rect 48495 27132 55146 27216
rect 48495 26964 48608 27132
rect 48776 26964 55146 27132
rect 48495 26880 55146 26964
rect 42280 26248 42963 26472
rect 42739 25339 42963 26248
rect -448 22078 783 22134
rect -448 22064 671 22078
rect -448 22008 -422 22064
rect -366 22022 671 22064
rect 727 22022 783 22078
rect -366 22008 783 22022
rect -448 21966 783 22008
rect 53312 20048 55146 26880
rect -11033 19961 -4087 20048
rect -11033 19793 -4368 19961
rect -4200 19793 -4087 19961
rect 48440 19962 55146 20048
rect -11033 19712 -4087 19793
rect 48440 19794 48552 19962
rect 48720 19794 55146 19962
rect 48440 19712 55146 19794
rect -11033 12880 -9199 19712
rect -224 18494 783 18550
rect -224 18480 671 18494
rect -224 18424 -196 18480
rect -140 18438 671 18480
rect 727 18438 783 18494
rect -140 18424 783 18438
rect -224 18382 783 18424
rect -280 14910 783 14966
rect -280 14896 671 14910
rect -280 14840 -195 14896
rect -139 14854 671 14896
rect 727 14854 783 14910
rect -139 14840 783 14854
rect -280 14798 783 14840
rect -4648 12880 -4592 12881
rect 53312 12880 55146 19712
rect -11033 12788 -4592 12880
rect -11033 12620 -4872 12788
rect -4704 12620 -4592 12788
rect 48552 12793 55146 12880
rect -11033 12544 -4592 12620
rect 48552 12625 48664 12793
rect 48832 12625 55146 12793
rect 48552 12544 55146 12625
rect -11033 5712 -9199 12544
rect -224 11326 783 11382
rect -224 11270 -202 11326
rect -146 11270 671 11326
rect 727 11270 783 11326
rect -224 11214 783 11270
rect -448 7799 -304 7800
rect -448 7798 -232 7799
rect -120 7798 -49 7799
rect -448 7742 783 7798
rect -448 7728 671 7742
rect -448 7672 -416 7728
rect -360 7686 671 7728
rect 727 7686 783 7742
rect -360 7672 783 7686
rect -448 7630 783 7672
rect 53312 5712 55146 12544
rect -11033 5623 -4032 5712
rect -11033 5455 -4312 5623
rect -4144 5455 -4032 5623
rect 48552 5627 55146 5712
rect -11033 5376 -4032 5455
rect 48552 5459 48664 5627
rect 48832 5459 55146 5627
rect 48552 5376 55146 5459
rect -11033 -4322 -9199 5376
rect -672 4158 783 4214
rect -672 4144 671 4158
rect -672 4088 -644 4144
rect -588 4102 671 4144
rect 727 4102 783 4158
rect -588 4088 783 4102
rect -672 4046 783 4088
rect -11033 -4326 -6226 -4322
rect 2139 -4326 2363 8
rect 3539 -1231 3763 239
rect 3192 -1348 4034 -1231
rect 3192 -1964 3306 -1348
rect 3924 -1964 4034 -1348
rect 3192 -2073 4034 -1964
rect 7739 -4326 7963 -1
rect 9139 -1231 9363 595
rect 8791 -1348 9633 -1231
rect 8791 -1964 8896 -1348
rect 9514 -1964 9633 -1348
rect 8791 -2073 9633 -1964
rect 13339 -4326 13563 -1
rect 14739 -1230 14963 1656
rect 14391 -1348 15233 -1230
rect 14391 -1964 14496 -1348
rect 15114 -1964 15233 -1348
rect 14391 -2072 15233 -1964
rect 18939 -4326 19163 19
rect 20339 -1038 20563 1816
rect 20338 -1230 20563 -1038
rect 20047 -1339 20889 -1230
rect 20047 -1955 20156 -1339
rect 20774 -1955 20889 -1339
rect 20047 -2072 20889 -1955
rect 24539 -4326 24763 -1
rect 25939 -1232 26163 938
rect 25595 -1339 26437 -1232
rect 25595 -1955 25706 -1339
rect 26324 -1955 26437 -1339
rect 25595 -2074 26437 -1955
rect 30139 -4326 30363 -1
rect 31538 -1230 31762 528
rect 31191 -1339 32033 -1230
rect 31191 -1955 31299 -1339
rect 31917 -1955 32033 -1339
rect 31191 -2072 32033 -1955
rect 35739 -4326 35963 0
rect 37139 -1230 37363 634
rect 36848 -1346 37690 -1230
rect 36848 -1962 36959 -1346
rect 37577 -1962 37690 -1346
rect 36848 -2072 37690 -1962
rect 41339 -4326 41563 0
rect 42739 -1230 42963 1189
rect 53312 686 55146 5376
rect 48440 595 55146 686
rect 48440 427 48577 595
rect 48745 427 55146 595
rect 48440 350 55146 427
rect 42448 -1342 43290 -1230
rect 42448 -1958 42560 -1342
rect 43178 -1958 43290 -1342
rect 42448 -2072 43290 -1958
rect 53312 -4324 55146 350
rect 51126 -4326 55146 -4324
rect -11033 -4872 55146 -4326
rect -11033 -6160 55143 -4872
rect -9904 -6161 -6226 -6160
rect 51126 -6163 55143 -6160
<< via3 >>
rect 3327 34775 3994 35401
rect 8907 34776 9574 35402
rect 20850 34776 21517 35402
rect 15400 32200 15512 32312
rect 25772 34778 26439 35404
rect 31321 34773 31988 35399
rect 36928 34774 37595 35400
rect 42168 34776 42785 35392
rect -4480 26956 -4312 27124
rect 2222 27018 2283 27078
rect 7822 27018 7883 27078
rect 13422 27018 13483 27078
rect 19022 27018 19083 27078
rect 24622 27018 24683 27078
rect 30222 27018 30283 27078
rect 48608 26964 48776 27132
rect 3617 23412 3678 23472
rect 9219 23406 9280 23466
rect 14818 23422 14879 23482
rect 20414 23403 20475 23463
rect 26020 23403 26081 23463
rect 31613 23400 31674 23460
rect 37211 23394 37272 23454
rect 42812 23411 42873 23471
rect -4368 19793 -4200 19961
rect 2222 19850 2283 19910
rect 7822 19850 7883 19910
rect 13422 19850 13483 19910
rect 19022 19850 19083 19910
rect 24622 19850 24683 19910
rect 30222 19850 30283 19910
rect 35822 19850 35883 19910
rect 41422 19850 41483 19910
rect 48552 19794 48720 19962
rect 3624 16223 3685 16283
rect 9220 16222 9281 16282
rect 14820 16223 14881 16283
rect 20420 16233 20481 16293
rect 26012 16222 26073 16282
rect 31624 16222 31685 16282
rect 37223 16230 37284 16290
rect 42817 16240 42878 16300
rect -3080 16139 -2968 16214
rect -4872 12620 -4704 12788
rect -2070 12662 -1942 12752
rect 2222 12682 2283 12742
rect 7822 12682 7883 12742
rect 13422 12682 13483 12742
rect 19022 12682 19083 12742
rect 24622 12682 24683 12742
rect 30222 12682 30283 12742
rect 35822 12682 35883 12742
rect 41422 12682 41483 12742
rect 48664 12625 48832 12793
rect 3621 9058 3682 9118
rect 9213 9058 9274 9118
rect 14819 9055 14880 9115
rect 20419 9063 20480 9123
rect 26019 9077 26080 9137
rect 31623 9055 31684 9115
rect 37217 9055 37278 9115
rect 42821 9074 42882 9134
rect -4312 5455 -4144 5623
rect 2222 5514 2283 5574
rect 7822 5514 7883 5574
rect 13422 5514 13483 5574
rect 19022 5514 19083 5574
rect 24622 5514 24683 5574
rect 30222 5514 30283 5574
rect 35822 5514 35883 5574
rect 41422 5514 41483 5574
rect 48664 5459 48832 5627
rect 3306 -1964 3924 -1348
rect 8896 -1964 9514 -1348
rect 14496 -1964 15114 -1348
rect 20156 -1955 20774 -1339
rect 25706 -1955 26324 -1339
rect 31299 -1955 31917 -1339
rect 36959 -1962 37577 -1346
rect 48577 427 48745 595
rect 42560 -1958 43178 -1342
<< metal4 >>
rect -7112 35404 51181 35992
rect -7112 35402 25772 35404
rect -7112 35401 8907 35402
rect -7112 34775 3327 35401
rect 3994 34776 8907 35401
rect 9574 34776 20850 35402
rect 21517 34778 25772 35402
rect 26439 35400 51181 35404
rect 26439 35399 36928 35400
rect 26439 34778 31321 35399
rect 21517 34776 31321 34778
rect 3994 34775 31321 34776
rect -7112 34773 31321 34775
rect 31988 34774 36928 35399
rect 37595 35392 51181 35400
rect 37595 34776 42168 35392
rect 42785 34776 51181 35392
rect 37595 34774 51181 34776
rect 31988 34773 51181 34774
rect -7112 34158 51181 34773
rect -7112 27217 -5278 34158
rect 15344 32312 15568 34158
rect 40008 34157 43890 34158
rect 15344 32200 15400 32312
rect 15512 32200 15568 32312
rect 15344 32144 15568 32200
rect -7112 26879 -5275 27217
rect -4281 27216 -2353 27217
rect 40083 27216 45741 27218
rect -4592 27132 48888 27216
rect -4592 27124 48608 27132
rect -4592 26956 -4480 27124
rect -4312 27078 48608 27124
rect -4312 27018 2222 27078
rect 2283 27018 7822 27078
rect 7883 27018 13422 27078
rect 13483 27018 19022 27078
rect 19083 27018 24622 27078
rect 24683 27018 30222 27078
rect 30283 27018 48608 27078
rect -4312 26964 48608 27018
rect 48776 26964 48888 27132
rect -4312 26956 48888 26964
rect -4592 26880 48888 26956
rect -4281 26879 -2353 26880
rect 40083 26879 45741 26880
rect -7112 23632 -5278 26879
rect 49336 23632 51181 34158
rect -7112 23482 51181 23632
rect -7112 23472 14818 23482
rect -7112 23412 3617 23472
rect 3678 23466 14818 23472
rect 3678 23412 9219 23466
rect -7112 23406 9219 23412
rect 9280 23422 14818 23466
rect 14879 23471 51181 23482
rect 14879 23463 42812 23471
rect 14879 23422 20414 23463
rect 9280 23406 20414 23422
rect -7112 23403 20414 23406
rect 20475 23403 26020 23463
rect 26081 23460 42812 23463
rect 26081 23403 31613 23460
rect -7112 23400 31613 23403
rect 31674 23454 42812 23460
rect 31674 23400 37211 23454
rect -7112 23394 37211 23400
rect 37272 23411 42812 23454
rect 42873 23411 51181 23471
rect 37272 23394 51181 23411
rect -7112 23296 51181 23394
rect -7112 16464 -5278 23296
rect 46898 23295 51181 23296
rect -4130 20049 -2379 20050
rect -4130 20048 46761 20049
rect -4480 19962 48833 20048
rect -4480 19961 48552 19962
rect -4480 19793 -4368 19961
rect -4200 19910 48552 19961
rect -4200 19850 2222 19910
rect 2283 19850 7822 19910
rect 7883 19850 13422 19910
rect 13483 19850 19022 19910
rect 19083 19850 24622 19910
rect 24683 19850 30222 19910
rect 30283 19850 35822 19910
rect 35883 19850 41422 19910
rect 41483 19850 48552 19910
rect -4200 19794 48552 19850
rect 48720 19794 48833 19962
rect -4200 19793 48833 19794
rect -4480 19713 48833 19793
rect -4480 19712 -2379 19713
rect 46732 19712 48833 19713
rect 49336 16465 51181 23295
rect 46762 16464 51181 16465
rect -7112 16300 51181 16464
rect -7112 16293 42817 16300
rect -7112 16283 20420 16293
rect -7112 16223 3624 16283
rect 3685 16282 14820 16283
rect 3685 16223 9220 16282
rect -7112 16222 9220 16223
rect 9281 16223 14820 16282
rect 14881 16233 20420 16283
rect 20481 16290 42817 16293
rect 20481 16282 37223 16290
rect 20481 16233 26012 16282
rect 14881 16223 26012 16233
rect 9281 16222 26012 16223
rect 26073 16222 31624 16282
rect 31685 16230 37223 16282
rect 37284 16240 42817 16290
rect 42878 16240 51181 16300
rect 37284 16230 51181 16240
rect 31685 16222 51181 16230
rect -7112 16214 51181 16222
rect -7112 16139 -3080 16214
rect -2968 16139 51181 16214
rect -7112 16128 51181 16139
rect -7112 9296 -5278 16128
rect -4648 12880 -4592 12881
rect -4130 12880 -2577 12881
rect -4985 12793 48944 12880
rect -4985 12788 48664 12793
rect -4985 12620 -4872 12788
rect -4704 12752 48664 12788
rect -4704 12662 -2070 12752
rect -1942 12742 48664 12752
rect -1942 12682 2222 12742
rect 2283 12682 7822 12742
rect 7883 12682 13422 12742
rect 13483 12682 19022 12742
rect 19083 12682 24622 12742
rect 24683 12682 30222 12742
rect 30283 12682 35822 12742
rect 35883 12682 41422 12742
rect 41483 12682 48664 12742
rect -1942 12662 48664 12682
rect -4704 12625 48664 12662
rect 48832 12625 48944 12793
rect -4704 12620 48944 12625
rect -4985 12544 48944 12620
rect -4130 12543 -2577 12544
rect 49336 9297 51181 16128
rect 46760 9296 51181 9297
rect -7112 9137 51181 9296
rect -7112 9123 26019 9137
rect -7112 9118 20419 9123
rect -7112 9058 3621 9118
rect 3682 9058 9213 9118
rect 9274 9115 20419 9118
rect 9274 9058 14819 9115
rect -7112 9055 14819 9058
rect 14880 9063 20419 9115
rect 20480 9077 26019 9123
rect 26080 9134 51181 9137
rect 26080 9115 42821 9134
rect 26080 9077 31623 9115
rect 20480 9063 31623 9077
rect 14880 9055 31623 9063
rect 31684 9055 37217 9115
rect 37278 9074 42821 9115
rect 42882 9074 51181 9134
rect 37278 9055 51181 9074
rect -7112 8960 51181 9055
rect -7112 2142 -5278 8960
rect -4131 5712 475 5714
rect -4424 5709 475 5712
rect 48552 5709 48944 5712
rect -4424 5627 48944 5709
rect -4424 5623 48664 5627
rect -4424 5455 -4312 5623
rect -4144 5574 48664 5623
rect -4144 5514 2222 5574
rect 2283 5514 7822 5574
rect 7883 5514 13422 5574
rect 13483 5514 19022 5574
rect 19083 5514 24622 5574
rect 24683 5514 30222 5574
rect 30283 5514 35822 5574
rect 35883 5514 41422 5574
rect 41483 5514 48664 5574
rect -4144 5459 48664 5514
rect 48832 5459 48944 5627
rect -4144 5455 48944 5459
rect -4424 5376 48944 5455
rect -1177 5373 48750 5376
rect 49336 2142 51181 8960
rect -7112 1806 -631 2142
rect -7112 -743 -5278 1806
rect 47012 1805 51181 2142
rect 47040 595 48867 686
rect 47040 427 48577 595
rect 48745 427 48867 595
rect 47040 350 48867 427
rect 49336 298 51181 1805
rect 49335 -743 51181 298
rect -7112 -1339 51181 -743
rect -7112 -1348 20156 -1339
rect -7112 -1964 3306 -1348
rect 3924 -1964 8896 -1348
rect 9514 -1964 14496 -1348
rect 15114 -1955 20156 -1348
rect 20774 -1955 25706 -1339
rect 26324 -1955 31299 -1339
rect 31917 -1342 51181 -1339
rect 31917 -1346 42560 -1342
rect 31917 -1955 36959 -1346
rect 15114 -1962 36959 -1955
rect 37577 -1958 42560 -1346
rect 43178 -1958 51181 -1342
rect 37577 -1962 51181 -1958
rect 15114 -1964 51181 -1962
rect -7112 -2577 51181 -1964
use 4MSB_weighted_binary  4MSB_weighted_binary_0
timestamp 1756789507
transform 1 0 36904 0 1 32033
box 2128 -3026 9800 1680
use 6MSB_MATRIX  6MSB_MATRIX_0
timestamp 1756722462
transform 1 0 951 0 1 -41314
box -1792 41313 46256 70567
use thermo_decoder  thermo_decoder_0
timestamp 1756615742
transform 0 1 14281 -1 0 33824
box 336 -337 3920 6440
use thermo_decoder  thermo_decoder_1
timestamp 1756615742
transform 1 0 -4592 0 1 11928
box 336 -337 3920 6440
<< labels >>
flabel metal4 -7112 34158 51165 35992 1 FreeSans 8000 0 0 0 VDD
port 15 n
flabel metal4 -7112 -2577 51176 -743 1 FreeSans 8000 0 0 0 VDD
port 15 n
flabel metal3 53312 -4872 55146 39636 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel metal3 -11033 -6160 55143 -4326 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel metal3 -11033 -6160 -9199 39636 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel metal3 -11033 37800 51109 39634 1 FreeSans 8000 0 0 0 VSS
port 16 n
rlabel metal3 49160 37802 55146 39636 1 VSS
flabel metal2 40435 41216 40595 41681 1 FreeSans 8000 0 0 0 X1
port 1 n
flabel metal2 34835 41180 34995 41645 1 FreeSans 8000 0 0 0 X2
port 2 n
flabel metal2 29236 41219 29396 41684 1 FreeSans 8000 0 0 0 X3
port 3 n
flabel metal2 23638 41164 23798 41629 1 FreeSans 8000 0 0 0 X4
port 4 n
flabel metal2 18090 41243 18250 41708 1 FreeSans 8000 0 0 0 X5
port 5 n
flabel metal2 7005 41227 7165 41692 1 FreeSans 8000 0 0 0 X7
port 7 n
flabel metal2 12548 41224 12708 41689 1 FreeSans 8000 0 0 0 X6
port 6 n
flabel metal2 1404 41184 1564 41649 1 FreeSans 8000 0 0 0 X10
port 10 n
flabel metal2 -3917 41201 -3757 41666 1 FreeSans 8000 0 0 0 X8
port 8 n
flabel metal2 -9795 41179 -9635 41644 1 FreeSans 8000 0 0 0 X9
port 9 n
flabel metal2 21678 41391 21831 41707 1 FreeSans 8000 0 0 0 CLK
port 11 n
flabel metal2 55664 34570 56056 34906 1 FreeSans 8000 0 0 0 OUTP
port 12 n
flabel metal2 60928 33929 61377 34266 1 FreeSans 8000 0 0 0 OUTN
port 13 n
flabel metal2 66248 33319 66697 33656 1 FreeSans 8000 0 0 0 VBIAS
port 14 n
flabel metal4 -7112 -2577 -5278 35992 1 FreeSans 8000 0 0 0 VDD
port 15 n
flabel metal4 49336 -2577 51181 35992 1 FreeSans 8000 0 0 0 VDD
port 15 n
<< end >>
