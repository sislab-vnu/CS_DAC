* NGSPICE file created from 4MSB_weighted_binary.ext - technology: gf180mcuD

.subckt CS_Switch_2x2 INP INN OUTP OUTN VBIAS VSS
X0 a_336_n248# VBIAS a_32_n20# VSS nfet_03v3 ad=0.2728p pd=1.905u as=0.1516p ps=1.64u w=0.22u l=0.28u
X1 OUTN INN a_32_n20# VSS nfet_03v3 ad=0.182p pd=1.8u as=0.102p ps=1u w=0.22u l=0.28u
X2 a_32_n20# INP OUTP VSS nfet_03v3 ad=0.102p pd=1u as=0.102p ps=1u w=0.22u l=0.28u
X3 OUTP VSS a_n246_n20# VSS nfet_03v3 ad=0.102p pd=1u as=50.6f ps=0.9u w=0.22u l=0.28u
X4 a_336_n248# VBIAS VSS VSS nfet_03v3 ad=0.2728p pd=1.905u as=0.132p ps=1.04u w=0.44u l=1.8u
X5 a_652_n20# VSS a_336_n248# VSS nfet_03v3 ad=50.6f pd=0.9u as=0.2728p ps=1.905u w=0.22u l=0.28u
X6 a_652_n248# VSS a_336_n248# VSS nfet_03v3 ad=0.1012p pd=1.34u as=0.2728p ps=1.905u w=0.44u l=0.28u
X7 VSS VSS a_n246_n248# VSS nfet_03v3 ad=0.132p pd=1.04u as=0.1012p ps=1.34u w=0.44u l=0.28u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
X0 VSS a_2304_115# Q VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1 VSS CLK a_36_151# VPW nfet_05v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2 Q a_2304_115# VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3 a_2304_115# a_2011_527# VSS VPW nfet_05v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4 a_1004_159# D a_836_159# VPW nfet_05v0 ad=0.207p pd=1.51u as=43.199997f ps=0.6u w=0.36u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_05v0 ad=0.1872p pd=1.4u as=53.999996f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_05v0 ad=0.1665p pd=1.285u as=0.1791p ps=1.355u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_05v0 ad=50.399998f pd=0.64u as=0.1665p ps=1.285u w=0.36u l=0.5u
X8 a_1376_115# a_1004_159# VDD VNW pfet_05v0 ad=0.1791p pd=1.355u as=0.1044p ps=0.94u w=0.36u l=0.5u
X9 VDD CLK a_36_151# VNW pfet_05v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X10 VDD a_2304_115# Q VNW pfet_05v0 ad=0.854p pd=3.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X11 VSS a_1376_115# a_1328_159# VPW nfet_05v0 ad=0.2637p pd=1.825u as=43.199997f ps=0.6u w=0.36u l=0.6u
X12 a_2011_527# a_448_472# a_1376_115# VPW nfet_05v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_05v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X14 Q a_2304_115# VDD VNW pfet_05v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X15 a_1376_115# a_1004_159# VSS VPW nfet_05v0 ad=93.59999f pd=0.88u as=0.2637p ps=1.825u w=0.36u l=0.6u
X16 VSS a_2304_115# a_2256_159# VPW nfet_05v0 ad=0.142p pd=1.14u as=43.199997f ps=0.6u w=0.36u l=0.6u
X17 a_836_159# a_36_151# VSS VPW nfet_05v0 ad=43.199997f pd=0.6u as=0.1584p ps=1.6u w=0.36u l=0.6u
X18 a_448_472# a_36_151# VSS VPW nfet_05v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X19 a_2256_159# a_36_151# a_2011_527# VPW nfet_05v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X20 a_880_527# a_448_472# VDD VNW pfet_05v0 ad=53.999996f pd=0.66u as=0.4554p ps=3.25u w=0.36u l=0.5u
X21 a_1348_527# a_36_151# a_1004_159# VNW pfet_05v0 ad=43.199997f pd=0.6u as=0.1872p ps=1.4u w=0.36u l=0.5u
X22 a_1328_159# a_448_472# a_1004_159# VPW nfet_05v0 ad=43.199997f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X23 VDD a_1376_115# a_1348_527# VNW pfet_05v0 ad=0.1044p pd=0.94u as=43.199997f ps=0.6u w=0.36u l=0.5u
X24 VDD a_2304_115# a_2296_527# VNW pfet_05v0 ad=0.23p pd=1.54u as=50.399998f ps=0.64u w=0.36u l=0.5u
X25 a_2304_115# a_2011_527# VDD VNW pfet_05v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt CS_Switch_8x2 INP INN OUTP OUTN VBIAS VSS
X0 a_784_1400# INP OUTP VSS nfet_03v3 ad=0.1306p pd=1.26u as=0.1328p ps=1.28u w=0.22u l=0.28u
X1 OUTP VSS a_450_1400# VSS nfet_03v3 ad=0.1328p pd=1.28u as=50.6f ps=0.9u w=0.22u l=0.28u
X2 OUTN INN a_784_1400# VSS nfet_03v3 ad=0.2106p pd=2.06u as=0.1306p ps=1.26u w=0.22u l=0.28u
X3 VSS VBIAS a_1348_1366# VSS nfet_03v3 ad=0.2026p pd=1.6u as=0.1357p ps=1.08u w=0.62u l=0.3u
X4 a_1348_1366# VBIAS a_784_1400# VSS nfet_03v3 ad=0.1357p pd=1.08u as=0.2248p ps=2.06u w=0.56u l=0.28u
X5 a_1712_1360# VSS VSS VSS nfet_03v3 ad=0.1426p pd=1.7u as=0.2026p ps=1.6u w=0.62u l=0.3u
.ends

.subckt CS_Switch_4x2 INP INN OUTP OUTN VBIAS VSS
X0 a_984_0# VSS a_812_0# VSS nfet_03v3 ad=0.1035p pd=1.36u as=0.1794p ps=1.525u w=0.45u l=0.28u
X1 a_42_240# INP OUTP VSS nfet_03v3 ad=0.102p pd=1u as=0.182p ps=1.8u w=0.22u l=0.28u
X2 a_812_0# VBIAS a_42_240# VSS nfet_03v3 ad=0.1794p pd=1.525u as=0.1516p ps=1.64u w=0.22u l=0.28u
X3 VSS VBIAS a_n110_0# VSS nfet_03v3 ad=0.2128p pd=1.78u as=0.1752p ps=1.48u w=0.45u l=1.8u
X4 a_n110_0# VSS a_n212_240# VSS nfet_03v3 ad=0.1752p pd=1.48u as=50.6f ps=0.9u w=0.22u l=0.28u
X5 a_42_240# VBIAS a_n110_0# VSS nfet_03v3 ad=0.1516p pd=1.64u as=0.1752p ps=1.48u w=0.22u l=0.28u
X6 a_984_240# VSS a_812_0# VSS nfet_03v3 ad=50.6f pd=0.9u as=0.1794p ps=1.525u w=0.22u l=0.28u
X7 OUTN INN a_42_240# VSS nfet_03v3 ad=0.182p pd=1.8u as=0.102p ps=1u w=0.22u l=0.28u
X8 a_n110_0# VSS a_n212_0# VSS nfet_03v3 ad=0.1752p pd=1.48u as=0.1035p ps=1.36u w=0.45u l=0.28u
X9 a_812_0# VBIAS VSS VSS nfet_03v3 ad=0.1794p pd=1.525u as=0.2128p ps=1.78u w=0.45u l=1.8u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
X0 Z a_36_68# VDD VNW pfet_05v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_05v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_05v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_05v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
X0 VDD I ZN VNW pfet_05v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_05v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_05v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
.ends

.subckt CS_Switch_1x1 INP INN OUTP OUTN VBIAS VSS
X0 a_668_n40# VSS a_440_n224# VSS nfet_03v3 ad=50.6f pd=0.9u as=0.1452p ps=1.465u w=0.22u l=0.28u
X1 a_668_n224# VSS a_440_n224# VSS nfet_03v3 ad=50.6f pd=0.9u as=0.1452p ps=1.465u w=0.22u l=0.28u
X2 a_440_n224# VBIAS a_56_n40# VSS nfet_03v3 ad=0.1452p pd=1.465u as=0.1516p ps=1.64u w=0.22u l=0.28u
X3 VSS VSS a_n228_n224# VSS nfet_03v3 ad=94.5f pd=0.99u as=50.6f ps=0.9u w=0.22u l=0.28u
X4 OUTN INN a_56_n40# VSS nfet_03v3 ad=0.182p pd=1.8u as=86.8f ps=0.92u w=0.22u l=0.28u
X5 a_440_n224# VBIAS VSS VSS nfet_03v3 ad=0.1452p pd=1.465u as=94.5f ps=0.99u w=0.22u l=2.2u
X6 a_56_n40# INP OUTP VSS nfet_03v3 ad=86.8f pd=0.92u as=0.1053p ps=1.03u w=0.22u l=0.28u
X7 OUTP VSS a_n228_n40# VSS nfet_03v3 ad=0.1053p pd=1.03u as=50.6f ps=0.9u w=0.22u l=0.28u
.ends

.subckt x4MSB_weighted_binary D1 D2 D3 D4 OUTP OUTN VBIAS CLK VDD VSS
XCS_Switch_2x2_1 CS_Switch_2x2_1/INP CS_Switch_2x2_1/INN OUTP OUTN VBIAS VSS CS_Switch_2x2
Xgf180mcu_fd_sc_mcu7t5v0__dffq_2_1 D1 CLK gf180mcu_fd_sc_mcu7t5v0__inv_2_1/I VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xgf180mcu_fd_sc_mcu7t5v0__dffq_2_0 D4 CLK gf180mcu_fd_sc_mcu7t5v0__inv_2_2/I VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xgf180mcu_fd_sc_mcu7t5v0__dffq_2_2 D2 CLK gf180mcu_fd_sc_mcu7t5v0__inv_2_0/I VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xgf180mcu_fd_sc_mcu7t5v0__dffq_2_3 D3 CLK gf180mcu_fd_sc_mcu7t5v0__inv_2_3/I VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_2
XCS_Switch_8x2_0 CS_Switch_8x2_0/INP CS_Switch_8x2_0/INN OUTP OUTN VBIAS VSS CS_Switch_8x2
XCS_Switch_4x2_0 CS_Switch_4x2_0/INP CS_Switch_4x2_0/INN OUTP OUTN VBIAS VSS CS_Switch_4x2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_0 gf180mcu_fd_sc_mcu7t5v0__buf_2_0/I CS_Switch_1x1_0/INN
+ VDD VDD gf180mcu_fd_sc_mcu7t5v0__buf_2_0/VPW VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xgf180mcu_fd_sc_mcu7t5v0__inv_2_0 gf180mcu_fd_sc_mcu7t5v0__inv_2_0/I gf180mcu_fd_sc_mcu7t5v0__buf_2_9/I
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xgf180mcu_fd_sc_mcu7t5v0__inv_2_1 gf180mcu_fd_sc_mcu7t5v0__inv_2_1/I gf180mcu_fd_sc_mcu7t5v0__buf_2_0/I
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_1 gf180mcu_fd_sc_mcu7t5v0__inv_2_2/I CS_Switch_8x2_0/INP
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xgf180mcu_fd_sc_mcu7t5v0__inv_2_2 gf180mcu_fd_sc_mcu7t5v0__inv_2_2/I gf180mcu_fd_sc_mcu7t5v0__buf_2_5/I
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xgf180mcu_fd_sc_mcu7t5v0__inv_2_3 gf180mcu_fd_sc_mcu7t5v0__inv_2_3/I gf180mcu_fd_sc_mcu7t5v0__buf_2_7/I
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_4 gf180mcu_fd_sc_mcu7t5v0__inv_2_3/I CS_Switch_4x2_0/INP
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_5 gf180mcu_fd_sc_mcu7t5v0__buf_2_5/I CS_Switch_8x2_0/INN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_6 gf180mcu_fd_sc_mcu7t5v0__inv_2_0/I CS_Switch_2x2_1/INP
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_7 gf180mcu_fd_sc_mcu7t5v0__buf_2_7/I CS_Switch_4x2_0/INN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_8 gf180mcu_fd_sc_mcu7t5v0__inv_2_1/I CS_Switch_1x1_0/INP
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xgf180mcu_fd_sc_mcu7t5v0__buf_2_9 gf180mcu_fd_sc_mcu7t5v0__buf_2_9/I CS_Switch_2x2_1/INN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XCS_Switch_1x1_0 CS_Switch_1x1_0/INP CS_Switch_1x1_0/INN OUTP OUTN VBIAS VSS CS_Switch_1x1
.ends

