magic
tech gf180mcuD
magscale 1 10
timestamp 1754386073
<< pwell >>
rect 1022 186 2056 266
rect 1022 124 1302 186
rect 1324 146 1404 186
rect 1304 124 1424 146
rect 1462 124 2056 186
rect 1022 -215 2056 124
rect 1022 -238 1424 -215
rect 1022 -278 1304 -238
rect 1324 -278 1404 -238
rect 1464 -278 2056 -215
rect 1022 -487 2056 -278
<< nmos >>
rect 1304 40 1424 100
rect 1584 -12 1640 100
rect 1732 -18 1792 106
rect 1304 -192 1424 -132
rect 1584 -192 1640 -80
rect 1732 -198 1792 -74
<< ndiff >>
rect 1324 178 1404 194
rect 1324 146 1340 178
rect 1304 130 1340 146
rect 1388 146 1404 178
rect 1388 130 1424 146
rect 1304 100 1424 130
rect 1686 100 1732 106
rect 1304 -6 1424 40
rect 1538 32 1584 100
rect 1516 -6 1584 32
rect 1324 -22 1404 -6
rect 1324 -70 1340 -22
rect 1388 -70 1404 -22
rect 1324 -86 1404 -70
rect 1480 -12 1584 -6
rect 1640 -12 1732 100
rect 1480 -22 1560 -12
rect 1480 -70 1496 -22
rect 1544 -70 1560 -22
rect 1480 -80 1560 -70
rect 1686 -18 1732 -12
rect 1792 26 1838 106
rect 1792 -6 1862 26
rect 1792 -18 1898 -6
rect 1818 -22 1898 -18
rect 1818 -70 1834 -22
rect 1882 -70 1898 -22
rect 1818 -74 1898 -70
rect 1686 -80 1732 -74
rect 1480 -86 1584 -80
rect 1304 -132 1424 -86
rect 1516 -124 1584 -86
rect 1538 -192 1584 -124
rect 1640 -192 1732 -80
rect 1304 -222 1424 -192
rect 1304 -238 1340 -222
rect 1324 -270 1340 -238
rect 1388 -238 1424 -222
rect 1686 -198 1732 -192
rect 1792 -86 1898 -74
rect 1792 -118 1862 -86
rect 1792 -198 1838 -118
rect 1388 -270 1404 -238
rect 1324 -286 1404 -270
<< ndiffc >>
rect 1340 130 1388 178
rect 1340 -70 1388 -22
rect 1496 -70 1544 -22
rect 1834 -70 1882 -22
rect 1340 -270 1388 -222
<< polysilicon >>
rect 1650 196 1730 212
rect 1650 162 1666 196
rect 1584 148 1666 162
rect 1714 162 1730 196
rect 1714 148 1792 162
rect 1178 100 1258 110
rect 1584 126 1792 148
rect 1584 100 1640 126
rect 1732 106 1792 126
rect 1178 94 1304 100
rect 1178 46 1194 94
rect 1242 46 1304 94
rect 1178 40 1304 46
rect 1424 40 1470 100
rect 1178 30 1258 40
rect 1584 -80 1640 -12
rect 1732 -74 1792 -18
rect 1178 -132 1258 -122
rect 1178 -138 1304 -132
rect 1178 -186 1194 -138
rect 1242 -186 1304 -138
rect 1178 -192 1304 -186
rect 1424 -192 1470 -132
rect 1178 -202 1258 -192
rect 1584 -238 1640 -192
rect 1732 -244 1792 -198
<< polycontact >>
rect 1666 148 1714 196
rect 1194 46 1242 94
rect 1194 -186 1242 -138
<< metal1 >>
rect 1652 203 1728 210
rect 1608 196 1769 203
rect 1326 186 1402 192
rect 1302 178 1462 186
rect 1302 130 1340 178
rect 1388 130 1462 178
rect 1608 148 1666 196
rect 1714 148 1769 196
rect 1608 137 1769 148
rect 1652 134 1728 137
rect 1302 124 1462 130
rect 1326 116 1402 124
rect 1180 104 1256 108
rect 1085 94 1256 104
rect 1085 46 1194 94
rect 1242 46 1256 94
rect 1085 38 1256 46
rect 1180 32 1256 38
rect 1326 -22 1402 -8
rect 1482 -22 1558 -8
rect 1326 -70 1340 -22
rect 1388 -70 1496 -22
rect 1544 -70 1558 -22
rect 1326 -84 1402 -70
rect 1482 -84 1558 -70
rect 1820 -22 1896 -8
rect 1820 -70 1834 -22
rect 1882 -70 1896 -22
rect 1820 -84 1896 -70
rect 1180 -131 1256 -124
rect 1085 -138 1256 -131
rect 1085 -186 1194 -138
rect 1242 -186 1256 -138
rect 1085 -197 1256 -186
rect 1180 -200 1256 -197
rect 1326 -216 1402 -208
rect 1304 -222 1456 -216
rect 1304 -270 1340 -222
rect 1388 -270 1456 -222
rect 1304 -278 1456 -270
rect 1326 -284 1402 -278
rect 1834 -332 1882 -84
rect 1176 -437 1966 -332
<< labels >>
flabel metal1 1608 137 1769 203 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 1400 -437 1966 -332 1 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional
flabel pwell 1196 -438 1308 -351 1 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
flabel metal1 1085 -197 1194 -131 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 1085 38 1194 104 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 1304 -278 1456 -216 1 FreeSans 400 0 0 0 OUTP
port 3 nsew signal bidirectional
flabel metal1 1302 124 1462 186 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
<< end >>
