VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CS_Switch_2x
  CLASS BLOCK ;
  FOREIGN CS_Switch_2x ;
  ORIGIN -3.435 -4.280 ;
  SIZE 7.970 BY 3.200 ;
  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.061600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.480 6.645 4.760 7.245 ;
    END
  END INP
  PIN INN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.061600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.620 6.650 5.900 7.250 ;
    END
  END INN
  PIN OUTP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.905 6.450 4.185 7.245 ;
        RECT 3.860 6.065 4.240 6.450 ;
    END
  END OUTP
  PIN OUTN
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.185 6.455 6.465 7.240 ;
        RECT 6.140 6.070 6.520 6.455 ;
    END
  END OUTN
  PIN VBIAS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 6.600 9.765 6.955 ;
    END
  END VBIAS
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 10.225 6.065 10.605 6.450 ;
        RECT 10.280 5.215 10.560 6.065 ;
        RECT 9.430 5.210 11.095 5.215 ;
        RECT 3.860 4.755 11.095 5.210 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.435 4.280 11.405 7.480 ;
    END
  END VPW
  OBS
      LAYER Metal1 ;
        RECT 5.000 6.070 5.380 6.455 ;
        RECT 6.825 6.070 7.205 6.455 ;
        RECT 5.040 5.810 5.320 6.070 ;
        RECT 6.880 5.810 7.160 6.070 ;
        RECT 5.035 5.530 7.160 5.810 ;
  END
END CS_Switch_2x
END LIBRARY

