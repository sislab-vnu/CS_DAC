magic
tech gf180mcuD
magscale 1 10
timestamp 1754908551
<< pwell >>
rect -377 631 825 1384
<< nmos >>
rect -204 1100 -144 1220
rect 126 1100 186 1220
rect 278 1100 338 1220
rect 608 1100 668 1220
rect -204 826 -144 950
rect 4 826 64 950
rect 130 832 186 944
rect 278 832 334 944
rect 400 826 460 950
rect 608 826 668 950
<< ndiff >>
rect -250 1100 -204 1220
rect -144 1183 126 1220
rect -144 1137 -32 1183
rect 14 1137 126 1183
rect -144 1100 126 1137
rect 186 1100 278 1220
rect 338 1183 608 1220
rect 338 1137 450 1183
rect 496 1137 608 1183
rect 338 1100 608 1137
rect 668 1100 714 1220
rect -250 826 -204 950
rect -144 924 -98 950
rect -42 924 4 950
rect -144 910 4 924
rect -144 864 -71 910
rect -25 864 4 910
rect -144 848 4 864
rect -144 826 -98 848
rect -42 826 4 848
rect 64 944 110 950
rect 210 944 254 1100
rect 354 944 400 950
rect 64 832 130 944
rect 186 832 278 944
rect 334 832 400 944
rect 64 826 110 832
rect 354 826 400 832
rect 460 924 506 950
rect 562 924 608 950
rect 460 910 608 924
rect 460 864 489 910
rect 535 864 608 910
rect 460 848 608 864
rect 460 826 506 848
rect 562 826 608 848
rect 668 826 714 950
<< ndiffc >>
rect -32 1137 14 1183
rect 450 1137 496 1183
rect -71 864 -25 910
rect 489 864 535 910
<< polysilicon >>
rect 116 1329 196 1346
rect 116 1283 133 1329
rect 179 1283 196 1329
rect 116 1266 196 1283
rect 268 1329 348 1346
rect 268 1283 285 1329
rect 331 1283 348 1329
rect 268 1266 348 1283
rect -204 1220 -144 1266
rect 126 1220 186 1266
rect 278 1220 338 1266
rect 608 1220 668 1266
rect -204 950 -144 1100
rect 126 1054 186 1100
rect -16 1033 64 1050
rect -16 987 1 1033
rect 47 1006 64 1033
rect 47 987 186 1006
rect -16 970 186 987
rect 4 950 64 970
rect 130 944 186 970
rect 278 1054 338 1100
rect 400 1033 480 1050
rect 400 1006 417 1033
rect 278 987 417 1006
rect 463 987 480 1033
rect 278 970 480 987
rect 278 944 334 970
rect 400 950 460 970
rect 608 950 668 1100
rect -204 780 -144 826
rect 4 780 64 826
rect 130 812 186 832
rect 278 812 334 832
rect -210 767 -138 780
rect 130 776 334 812
rect 400 780 460 826
rect 608 780 668 826
rect -210 721 -197 767
rect -151 721 -138 767
rect -210 708 -138 721
rect 602 767 674 780
rect 602 721 615 767
rect 661 721 674 767
rect 602 708 674 721
<< polycontact >>
rect 133 1283 179 1329
rect 285 1283 331 1329
rect 1 987 47 1033
rect 417 987 463 1033
rect -197 721 -151 767
rect 615 721 661 767
<< metal1 >>
rect 118 1329 194 1344
rect 118 1283 133 1329
rect 179 1283 194 1329
rect 118 1268 194 1283
rect 270 1329 346 1344
rect 270 1283 285 1329
rect 331 1283 346 1329
rect 270 1268 346 1283
rect -47 1183 29 1198
rect -47 1137 -32 1183
rect 14 1137 29 1183
rect -47 1122 29 1137
rect 435 1183 511 1198
rect 435 1137 450 1183
rect 496 1137 511 1183
rect 435 1122 511 1137
rect -14 1033 62 1048
rect -14 987 1 1033
rect 47 987 62 1033
rect -14 972 62 987
rect 402 1033 478 1048
rect 402 987 417 1033
rect 463 987 478 1033
rect 402 972 478 987
rect -71 910 -25 921
rect -71 810 -25 864
rect 489 910 535 921
rect 489 810 535 864
rect -294 767 756 810
rect -294 721 -197 767
rect -151 721 615 767
rect 661 721 756 767
rect -294 690 756 721
<< labels >>
flabel metal1 118 1268 194 1344 1 FreeSans 400 0 0 0 INP
port 1 n
flabel metal1 270 1268 346 1344 1 FreeSans 400 0 0 0 INN
port 2 n
flabel metal1 -47 1122 29 1198 1 FreeSans 400 0 0 0 OUTP
port 3 n
flabel metal1 435 1122 511 1198 1 FreeSans 400 0 0 0 OUTN
port 4 n
flabel metal1 -14 972 62 1048 1 FreeSans 400 0 0 0 VBIAS
port 5 n
flabel metal1 402 972 478 1048 1 FreeSans 400 0 0 0 VBIAS
port 6 n
flabel metal1 -151 690 615 810 1 FreeSans 400 0 0 0 VSS
port 7 n
flabel pwell -327 688 -224 814 1 FreeSans 400 0 0 0 VPW
port 8 n
<< end >>
