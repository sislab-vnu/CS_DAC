magic
tech gf180mcuD
magscale 1 10
timestamp 1755857852
<< pwell >>
rect 31079 8826 31192 8882
<< metal1 >>
rect 11159 35544 11979 35850
rect 11159 35293 11420 35544
rect 11741 35293 11979 35544
rect 11159 35023 11979 35293
rect 11424 26544 11760 35023
rect 25536 26742 25872 26880
rect 25536 26686 25676 26742
rect 25732 26686 25872 26742
rect 25536 26544 25872 26686
rect 38917 26600 39256 26656
rect 33880 26544 39256 26600
rect 11480 25928 11704 26544
rect -952 25592 11704 25928
rect -952 20425 -615 25592
rect 9799 25370 10404 25371
rect 13247 25370 14416 25372
rect 25592 25370 25816 26544
rect 33880 26468 39032 26544
rect 33879 26432 39032 26468
rect 39144 26432 39256 26544
rect 33879 26320 39256 26432
rect 33879 26039 34162 26320
rect 41269 26264 41609 26377
rect 41269 26152 41384 26264
rect 41496 26152 41609 26264
rect 41269 26041 41609 26152
rect 41273 26040 41608 26041
rect -392 25034 29848 25370
rect -392 25033 11497 25034
rect 12181 25033 29848 25034
rect -316 24043 -221 25033
rect -133 24829 -37 24925
rect -133 24774 -112 24829
rect -56 24774 -37 24829
rect -133 24293 -37 24774
rect -317 23882 -221 24043
rect -132 24041 -37 24293
rect 8287 24152 8395 25033
rect 8287 24085 8300 24152
rect 8381 24085 8395 24152
rect 8287 24071 8395 24085
rect 18009 24128 18091 25033
rect 18009 24076 18021 24128
rect 18079 24076 18091 24128
rect 28146 24178 28216 25033
rect 28146 24122 28151 24178
rect 28207 24122 28216 24178
rect 28146 24108 28216 24122
rect -133 23969 -37 24041
rect -317 23614 -222 23882
rect -133 23788 -38 23969
rect -133 23707 -37 23788
rect -318 23420 -222 23614
rect -318 23147 -223 23420
rect -132 23261 -37 23707
rect 30681 23688 34107 24024
rect 30943 23687 31522 23688
rect 28147 23572 28213 23586
rect 18014 23527 18085 23539
rect -132 23166 309 23261
rect 8287 23236 8395 23300
rect -132 23165 -37 23166
rect -318 22991 -221 23147
rect 8287 23168 8307 23236
rect 8379 23168 8395 23236
rect -316 22753 -221 22991
rect -317 22524 -221 22753
rect 8287 22819 8395 23168
rect 8589 23243 9036 23274
rect 8589 23169 8680 23243
rect 8793 23169 9036 23243
rect 8589 23154 9036 23169
rect 13825 23240 15130 23274
rect 13825 23184 13888 23240
rect 13944 23184 15130 23240
rect 13825 23154 15130 23184
rect 8287 22721 9191 22819
rect 18014 22800 18085 23471
rect 28147 23520 28155 23572
rect 28208 23520 28213 23572
rect 18192 23240 18753 23274
rect 18192 23184 18283 23240
rect 18339 23184 18753 23240
rect 18192 23154 18753 23184
rect 23438 23240 24803 23274
rect 23438 23184 23493 23240
rect 23549 23184 24803 23240
rect 23438 23154 24803 23184
rect 28147 22852 28213 23520
rect 29296 23154 29448 23274
rect 18014 22729 18820 22800
rect 28147 22786 28508 22852
rect 8287 22720 8395 22721
rect -317 22225 -222 22524
rect 11045 22465 11946 22491
rect 11045 22389 11761 22465
rect 11874 22389 11946 22465
rect 11045 22369 11946 22389
rect 15764 22456 16758 22490
rect 15764 22400 16605 22456
rect 16661 22400 16758 22456
rect 15764 22368 16758 22400
rect 20732 22456 21585 22490
rect 20732 22400 21421 22456
rect 21477 22400 21585 22456
rect 20732 22370 21585 22400
rect 25777 22456 26400 22490
rect 25777 22400 26292 22456
rect 26348 22400 26400 22456
rect 25777 22370 26400 22400
rect 30382 22456 31263 22490
rect 30382 22400 31111 22456
rect 31167 22400 31263 22456
rect 30382 22370 31263 22400
rect -317 22130 306 22225
rect -952 20350 307 20425
rect -952 15780 -615 20350
rect 6040 19995 6311 20115
rect 6042 17195 6313 17315
rect -952 15721 287 15780
rect -952 10248 -615 15721
rect 5995 14395 6266 14515
rect 6832 13374 7056 13403
rect 6832 13305 6885 13374
rect 7001 13305 7056 13374
rect 6832 13283 7056 13305
rect 6046 11595 6317 11715
rect -952 10180 297 10248
rect -952 4582 -615 10180
rect 27833 9733 28055 9762
rect 27833 9663 27888 9733
rect 28000 9663 28055 9733
rect 27833 9634 28055 9663
rect 6046 8795 6317 8915
rect 27831 6939 28053 6967
rect 27831 6869 27887 6939
rect 27999 6869 28053 6939
rect 27831 6832 28053 6869
rect 6047 5995 6318 6115
rect -952 4521 330 4582
rect -952 2800 -615 4521
rect 6052 3195 6323 3315
rect 6043 395 6314 515
<< via1 >>
rect 11420 35293 11741 35544
rect 25676 26686 25732 26742
rect 39032 26432 39144 26544
rect 35783 26137 35896 26199
rect 41384 26152 41496 26264
rect 37139 25335 37230 25411
rect 35784 25176 35897 25238
rect -112 24774 -56 24829
rect 8300 24085 8381 24152
rect 18021 24076 18079 24128
rect 37137 24378 37228 24454
rect 35784 24221 35896 24283
rect 28151 24122 28207 24178
rect 18014 23471 18085 23527
rect 470 23133 526 23187
rect 8307 23168 8379 23236
rect 8680 23169 8793 23243
rect 13888 23184 13944 23240
rect 391 22657 504 22733
rect 9350 22790 9409 22850
rect 10361 22794 10415 22848
rect 15127 22763 15182 22816
rect 28155 23520 28208 23572
rect 18283 23184 18339 23240
rect 23493 23184 23549 23240
rect 37140 23426 37220 23495
rect 28442 23177 28542 23245
rect 35784 23238 35896 23300
rect 18982 22794 19043 22850
rect 24918 22793 24979 22852
rect 28671 22793 28732 22850
rect 29788 22792 29852 22852
rect 3881 22614 3971 22672
rect 11761 22389 11874 22465
rect 16605 22400 16661 22456
rect 21421 22400 21477 22456
rect 26292 22400 26348 22456
rect 31111 22400 31167 22456
rect 37137 22449 37216 22518
rect 4090 22229 4144 22282
rect 3865 22172 3920 22224
rect 2184 21703 2296 21777
rect 6887 21698 7001 21776
rect 11760 21700 11873 21782
rect 16593 21710 16683 21769
rect 21412 21709 21490 21773
rect 26264 21706 26375 21776
rect 31080 21714 31193 21771
rect 37146 21707 37224 21773
rect 244 21380 302 21434
rect 470 21325 525 21377
rect 392 20849 505 20925
rect 3864 20871 3976 20940
rect 8678 20855 8793 20940
rect 13889 20866 14003 20934
rect 18268 20864 18348 20943
rect 23462 20862 23576 20944
rect 27887 20864 28000 20937
rect 33039 20874 33155 20938
rect 35784 20869 35896 20928
rect 2184 20019 2296 20085
rect 6888 20014 7000 20091
rect 11760 20016 11872 20098
rect 16583 20022 16673 20081
rect 21409 20021 21486 20085
rect 26277 20017 26366 20089
rect 31079 20020 31192 20077
rect 37145 20023 37223 20089
rect 2184 18907 2296 18973
rect 6888 18901 7000 18976
rect 11760 18904 11872 18986
rect 16593 18910 16665 18969
rect 21404 18914 21481 18978
rect 26281 18903 26370 18975
rect 31080 18911 31192 18969
rect 37151 18909 37227 18978
rect 392 18005 505 18072
rect 3863 18059 3977 18136
rect 8680 18055 8792 18139
rect 13888 18070 14002 18138
rect 18269 18065 18349 18144
rect 23464 18068 23575 18143
rect 27889 18066 28002 18139
rect 33038 18053 33154 18117
rect 35784 18068 35896 18127
rect 454 17621 510 17673
rect 231 17561 284 17616
rect 2184 17214 2296 17300
rect 6888 17221 7000 17291
rect 11761 17212 11872 17282
rect 16599 17219 16671 17278
rect 21407 17212 21487 17285
rect 26270 17214 26369 17285
rect 31080 17221 31192 17279
rect 37143 17220 37219 17289
rect 2184 16117 2296 16181
rect 6887 16104 7000 16173
rect 11762 16110 11873 16180
rect 16588 16114 16667 16175
rect 21411 16108 21491 16181
rect 26271 16105 26370 16176
rect 31080 16115 31192 16171
rect 37144 16111 37218 16175
rect 450 15724 505 15779
rect 378 15254 513 15321
rect 3863 15255 3977 15332
rect 8679 15249 8791 15343
rect 13887 15263 14008 15338
rect 18267 15261 18351 15336
rect 23462 15258 23577 15324
rect 27888 15263 28000 15334
rect 33040 15269 33152 15339
rect 35784 15274 35896 15333
rect 2184 14425 2296 14495
rect 6888 14420 7001 14489
rect 11760 14418 11873 14494
rect 16592 14417 16671 14478
rect 21397 14410 21484 14481
rect 26265 14414 26371 14483
rect 31080 14423 31192 14479
rect 37150 14425 37224 14489
rect 2184 13310 2296 13383
rect 6885 13305 7001 13374
rect 11760 13308 11873 13384
rect 16594 13308 16668 13372
rect 21406 13305 21493 13376
rect 26267 13311 26373 13380
rect 31080 13310 31192 13370
rect 37148 13308 37226 13376
rect 3864 12464 3977 12535
rect 396 12402 501 12463
rect 8681 12455 8793 12549
rect 13885 12460 14006 12535
rect 18268 12455 18352 12530
rect 23462 12460 23577 12526
rect 27889 12456 28001 12527
rect 33040 12465 33152 12535
rect 35784 12465 35896 12524
rect 450 11987 507 12043
rect 2184 11616 2296 11700
rect 6886 11615 7002 11684
rect 11760 11611 11872 11686
rect 16601 11617 16675 11681
rect 21397 11610 21483 11686
rect 26278 11611 26367 11687
rect 31080 11625 31192 11685
rect 37146 11618 37224 11686
rect 2184 10503 2296 10581
rect 6887 10505 7001 10576
rect 11760 10508 11872 10583
rect 16593 10512 16669 10574
rect 21402 10500 21488 10576
rect 26277 10506 26366 10582
rect 31080 10518 31193 10573
rect 37137 10506 37219 10579
rect 461 10123 516 10178
rect 368 9654 474 9719
rect 3863 9670 3976 9741
rect 8680 9647 8794 9730
rect 13887 9663 14004 9735
rect 18265 9655 18353 9735
rect 23463 9663 23578 9726
rect 27888 9663 28000 9733
rect 33031 9666 33143 9732
rect 35784 9674 35896 9732
rect 347 9217 404 9274
rect 2184 8813 2296 8893
rect 6886 8814 7000 8885
rect 11760 8811 11872 8889
rect 16598 8816 16674 8878
rect 21397 8811 21484 8885
rect 26265 8811 26364 8886
rect 31079 8826 31192 8882
rect 37142 8812 37224 8885
rect 2184 7714 2296 7784
rect 6888 7708 7000 7773
rect 11760 7703 11872 7781
rect 16589 7706 16670 7772
rect 21404 7705 21491 7779
rect 26273 7708 26372 7783
rect 31079 7716 31192 7772
rect 37144 7711 37228 7779
rect 390 6805 505 6874
rect 3863 6854 3977 6935
rect 8679 6849 8791 6928
rect 13886 6866 14003 6938
rect 18263 6876 18351 6956
rect 23462 6865 23577 6928
rect 27887 6869 27999 6939
rect 33041 6864 33153 6930
rect 35784 6863 35896 6921
rect 334 6421 389 6473
rect 554 6416 618 6479
rect 2184 6012 2296 6088
rect 6888 6016 7000 6081
rect 11761 6016 11874 6089
rect 16593 6016 16674 6082
rect 21400 6011 21485 6083
rect 26275 6010 26367 6090
rect 31080 6026 31193 6082
rect 37140 6015 37224 6083
rect 2184 4910 2296 4984
rect 6888 4903 7001 4974
rect 11759 4907 11872 4980
rect 16589 4906 16672 4976
rect 21408 4902 21493 4974
rect 26281 4900 26373 4980
rect 31080 4921 31192 4977
rect 37140 4910 37228 4976
rect 557 4523 611 4577
rect 390 4062 507 4141
rect 3863 4058 3977 4139
rect 8680 4052 8793 4129
rect 13887 4060 14000 4135
rect 18267 4066 18360 4141
rect 23460 4056 23576 4127
rect 27887 4050 28001 4123
rect 33030 4072 33139 4136
rect 35783 4074 35896 4130
rect 333 3620 388 3674
rect 2184 3214 2296 3293
rect 6888 3217 7001 3288
rect 11757 3209 11875 3284
rect 16594 3218 16677 3288
rect 21401 3212 21486 3283
rect 26264 3210 26360 3290
rect 31080 3222 31192 3278
rect 37137 3219 37225 3285
rect 2184 2104 2296 2172
rect 6887 2104 7001 2173
rect 11758 2106 11876 2181
rect 16595 2104 16675 2177
rect 21403 2103 21488 2174
rect 26276 2099 26372 2179
rect 31079 2117 31193 2178
rect 3864 1265 3976 1332
rect 8679 1257 8792 1334
rect 13872 1255 14002 1328
rect 18262 1260 18355 1335
rect 23462 1271 23578 1342
rect 27887 1257 28001 1330
rect 33043 1265 33152 1329
rect 2184 416 2296 489
rect 6887 418 7001 487
rect 11760 410 11872 487
rect 16588 412 16668 485
rect 21402 408 21481 480
rect 26275 406 26363 483
rect 31079 421 31193 482
<< metal2 >>
rect 8112 35100 8932 35927
rect 11159 35544 11979 35850
rect 11159 35293 11420 35544
rect 11741 35293 11979 35544
rect 8344 26544 8680 35100
rect 11159 35023 11979 35293
rect 21602 35265 22422 36092
rect 25299 35318 26119 36145
rect 21840 26544 22176 35265
rect 25536 26742 25872 35318
rect 29980 35246 30800 36073
rect 31704 35276 32524 36103
rect 33185 35283 34005 36110
rect 25536 26686 25676 26742
rect 25732 26686 25872 26742
rect 25536 26544 25872 26686
rect 30184 26544 30520 35246
rect 31920 26544 32256 35276
rect 33432 26544 33768 35283
rect 34937 35280 35757 36107
rect 35168 26880 35504 35280
rect 38668 35091 39488 35918
rect 8400 26376 8625 26544
rect -1344 26371 8625 26376
rect -1344 26040 8624 26371
rect -1344 21444 -1007 26040
rect 11535 24977 12172 24978
rect 21896 24977 22120 26544
rect -168 24829 30072 24977
rect -168 24774 -112 24829
rect -56 24774 30072 24829
rect -168 24641 30072 24774
rect -168 24640 13276 24641
rect 14319 24640 30072 24641
rect 453 24380 548 24499
rect 453 24324 472 24380
rect 530 24324 548 24380
rect 453 23187 548 24324
rect 453 23133 470 23187
rect 526 23133 548 23187
rect 453 23121 548 23133
rect 336 22733 562 22762
rect 336 22657 391 22733
rect 504 22657 562 22733
rect 336 22628 562 22657
rect 3836 22672 4021 22707
rect 3836 22614 3881 22672
rect 3971 22614 4021 22672
rect 3836 22586 4021 22614
rect 4080 22292 4152 24640
rect 8287 24152 8395 24160
rect 8287 24085 8300 24152
rect 8381 24085 8395 24152
rect 8287 23258 8395 24085
rect 8272 23236 8403 23258
rect 8272 23168 8307 23236
rect 8379 23168 8403 23236
rect 8272 23148 8403 23168
rect 8624 23243 8847 23275
rect 8624 23169 8680 23243
rect 8793 23169 8847 23243
rect 8624 23154 8847 23169
rect 9342 22857 9414 24640
rect 13878 23240 13954 23250
rect 13878 23184 13888 23240
rect 13944 23184 13954 23240
rect 13878 23174 13954 23184
rect 9327 22850 9428 22857
rect 9327 22790 9350 22850
rect 9409 22790 9428 22850
rect 9327 22785 9428 22790
rect 10348 22850 10428 22860
rect 10348 22792 10358 22850
rect 10418 22792 10428 22850
rect 15121 22828 15185 24640
rect 18014 24128 18085 24140
rect 18014 24076 18021 24128
rect 18079 24076 18085 24128
rect 18014 23541 18085 24076
rect 17999 23527 18095 23541
rect 17999 23471 18014 23527
rect 18085 23471 18095 23527
rect 17999 23462 18095 23471
rect 18273 23240 18349 23250
rect 18273 23184 18283 23240
rect 18339 23184 18349 23240
rect 18273 23174 18349 23184
rect 18976 22856 19048 24640
rect 23483 23240 23559 23250
rect 23483 23184 23493 23240
rect 23549 23184 23559 23240
rect 23483 23174 23559 23184
rect 24912 22860 24984 24640
rect 28137 24178 28222 24185
rect 28137 24124 28151 24178
rect 28147 24122 28151 24124
rect 28207 24124 28222 24178
rect 28207 24122 28213 24124
rect 28147 23582 28213 24122
rect 28133 23572 28228 23582
rect 28133 23520 28155 23572
rect 28208 23520 28228 23572
rect 28133 23509 28228 23520
rect 27833 23261 28448 23262
rect 27833 23260 28553 23261
rect 27833 23251 28555 23260
rect 27833 23179 27862 23251
rect 28000 23245 28555 23251
rect 28000 23179 28442 23245
rect 27833 23177 28442 23179
rect 28542 23177 28555 23245
rect 27833 23167 28555 23177
rect 27938 23166 28555 23167
rect 28427 23164 28555 23166
rect 18968 22850 19057 22856
rect 10348 22782 10428 22792
rect 15114 22816 15195 22828
rect 15114 22763 15127 22816
rect 15182 22763 15195 22816
rect 18968 22794 18982 22850
rect 19043 22794 19057 22850
rect 18968 22788 19057 22794
rect 24905 22852 24993 22860
rect 28662 22855 28734 24640
rect 30240 23576 30464 26544
rect 31976 25978 32200 26544
rect 31976 23968 32201 25978
rect 33488 24920 33712 26544
rect 35224 25571 35448 26880
rect 38920 26544 39256 35091
rect 51734 27384 52331 27523
rect 40768 27047 52331 27384
rect 40768 27016 41104 27047
rect 40767 27015 41104 27016
rect 40767 26709 41103 27015
rect 51734 26958 52331 27047
rect 38920 26432 39032 26544
rect 39144 26432 39256 26544
rect 38920 26320 39256 26432
rect 40766 26680 41103 26709
rect 40766 26373 41102 26680
rect 41269 26264 41609 26377
rect 35728 26199 35952 26214
rect 35728 26137 35783 26199
rect 35896 26137 35952 26199
rect 41269 26161 41384 26264
rect 35728 26113 35952 26137
rect 41268 26152 41384 26161
rect 41496 26152 41609 26264
rect 41268 25864 41609 26152
rect 52349 25864 52946 25989
rect 41268 25527 52946 25864
rect 41307 25526 52946 25527
rect 37095 25411 37276 25429
rect 52349 25424 52946 25526
rect 37095 25335 37139 25411
rect 37230 25335 37276 25411
rect 37095 25320 37276 25335
rect 35750 25238 35928 25254
rect 35750 25176 35784 25238
rect 35897 25176 35928 25238
rect 35750 25154 35928 25176
rect 33488 24696 35319 24920
rect 37085 24454 37283 24467
rect 37085 24378 37137 24454
rect 37228 24378 37283 24454
rect 37085 24368 37283 24378
rect 35748 24283 35926 24295
rect 35748 24221 35784 24283
rect 35896 24221 35926 24283
rect 35748 24195 35926 24221
rect 31976 23744 35336 23968
rect 30240 23352 35432 23576
rect 37085 23495 37283 23510
rect 37085 23426 37140 23495
rect 37220 23426 37283 23495
rect 37085 23411 37283 23426
rect 30846 23349 31575 23352
rect 24905 22793 24918 22852
rect 24979 22793 24993 22852
rect 24905 22785 24993 22793
rect 28648 22850 28750 22855
rect 28648 22793 28671 22850
rect 28732 22793 28750 22850
rect 28648 22784 28750 22793
rect 29778 22852 29862 22862
rect 29778 22792 29788 22852
rect 29852 22792 29862 22852
rect 29778 22782 29862 22792
rect 15114 22752 15195 22763
rect 35208 22728 35432 23352
rect 35739 23300 35940 23321
rect 35739 23238 35784 23300
rect 35896 23238 35940 23300
rect 35739 23218 35940 23238
rect 37101 22518 37264 22537
rect 11727 22465 11904 22491
rect 11727 22389 11761 22465
rect 11874 22389 11904 22465
rect 16595 22456 16671 22466
rect 16595 22400 16605 22456
rect 16661 22400 16671 22456
rect 16595 22390 16671 22400
rect 21411 22456 21487 22466
rect 21411 22400 21421 22456
rect 21477 22400 21487 22456
rect 21411 22390 21487 22400
rect 26282 22456 26358 22466
rect 26282 22400 26292 22456
rect 26348 22400 26358 22456
rect 26282 22390 26358 22400
rect 31101 22456 31177 22466
rect 31101 22400 31111 22456
rect 31167 22400 31177 22456
rect 37101 22449 37137 22518
rect 37216 22449 37264 22518
rect 37101 22436 37264 22449
rect 31101 22390 31177 22400
rect 11727 22369 11904 22389
rect 4067 22282 4162 22292
rect 3851 22226 3934 22237
rect 3851 22170 3862 22226
rect 3923 22170 3934 22226
rect 4067 22229 4090 22282
rect 4144 22229 4162 22282
rect 4067 22213 4162 22229
rect 3851 22159 3934 22170
rect 2128 21777 2352 21803
rect 2128 21703 2184 21777
rect 2296 21703 2352 21777
rect 2128 21683 2352 21703
rect 6832 21776 7056 21803
rect 6832 21698 6887 21776
rect 7001 21698 7056 21776
rect 6832 21683 7056 21698
rect 11704 21782 11928 21803
rect 11704 21700 11760 21782
rect 11873 21700 11928 21782
rect 11704 21683 11928 21700
rect 16520 21769 16744 21803
rect 16520 21710 16593 21769
rect 16683 21710 16744 21769
rect 16520 21683 16744 21710
rect 21358 21773 21543 21792
rect 21358 21709 21412 21773
rect 21490 21709 21543 21773
rect 21358 21696 21543 21709
rect 26222 21776 26412 21792
rect 26222 21706 26264 21776
rect 26375 21706 26412 21776
rect 26222 21687 26412 21706
rect 31024 21771 31248 21792
rect 31024 21714 31080 21771
rect 31193 21714 31248 21771
rect 31024 21691 31248 21714
rect 37107 21773 37270 21793
rect 37107 21707 37146 21773
rect 37224 21707 37270 21773
rect 37107 21692 37270 21707
rect 230 21444 320 21449
rect -1344 21434 320 21444
rect -1344 21380 244 21434
rect 302 21380 320 21434
rect -1344 21376 320 21380
rect -1344 17545 -1007 21376
rect 230 21372 320 21376
rect 457 21380 538 21390
rect 457 21323 467 21380
rect 528 21323 538 21380
rect 457 21313 538 21323
rect 335 20925 559 20947
rect 335 20849 392 20925
rect 505 20849 559 20925
rect 335 20829 559 20849
rect 3808 20940 4034 20970
rect 3808 20871 3864 20940
rect 3976 20871 4034 20940
rect 3808 20844 4034 20871
rect 8623 20940 8848 20987
rect 8623 20855 8678 20940
rect 8793 20855 8848 20940
rect 8623 20822 8848 20855
rect 13856 20934 14035 20958
rect 13856 20866 13889 20934
rect 14003 20866 14035 20934
rect 13856 20835 14035 20866
rect 18231 20943 18383 20974
rect 18231 20864 18268 20943
rect 18348 20864 18383 20943
rect 18231 20834 18383 20864
rect 23408 20944 23632 20973
rect 23408 20862 23462 20944
rect 23576 20862 23632 20944
rect 23408 20832 23632 20862
rect 27831 20937 28057 20949
rect 27831 20864 27887 20937
rect 28000 20864 28057 20937
rect 27831 20833 28057 20864
rect 32984 20938 33208 20974
rect 32984 20874 33039 20938
rect 33155 20874 33208 20938
rect 32984 20848 33208 20874
rect 35736 20928 35937 20948
rect 35736 20869 35784 20928
rect 35896 20869 35937 20928
rect 35736 20845 35937 20869
rect 2128 20085 2352 20115
rect 2128 20019 2184 20085
rect 2296 20019 2352 20085
rect 2128 19995 2352 20019
rect 6832 20091 7057 20115
rect 6832 20014 6888 20091
rect 7000 20014 7057 20091
rect 6832 19995 7057 20014
rect 11704 20098 11928 20115
rect 11704 20016 11760 20098
rect 11872 20016 11928 20098
rect 11704 19995 11928 20016
rect 16540 20081 16720 20096
rect 16540 20022 16583 20081
rect 16673 20022 16720 20081
rect 16540 20004 16720 20022
rect 21355 20085 21540 20098
rect 21355 20021 21409 20085
rect 21486 20021 21540 20085
rect 21355 20006 21540 20021
rect 26228 20089 26418 20104
rect 26228 20017 26277 20089
rect 26366 20017 26418 20089
rect 26228 19999 26418 20017
rect 31023 20077 31248 20097
rect 31023 20020 31079 20077
rect 31192 20020 31248 20077
rect 31023 20003 31248 20020
rect 37092 20089 37277 20108
rect 37092 20023 37145 20089
rect 37223 20023 37277 20089
rect 37092 20006 37277 20023
rect 2128 18973 2352 19003
rect 2128 18907 2184 18973
rect 2296 18907 2352 18973
rect 2128 18883 2352 18907
rect 6832 18976 7056 19002
rect 6832 18901 6888 18976
rect 7000 18901 7056 18976
rect 6832 18883 7056 18901
rect 11704 18986 11928 19002
rect 11704 18904 11760 18986
rect 11872 18904 11928 18986
rect 11704 18883 11928 18904
rect 16540 18969 16720 18988
rect 16540 18910 16593 18969
rect 16665 18910 16720 18969
rect 16540 18896 16720 18910
rect 21371 18978 21516 18995
rect 21371 18914 21404 18978
rect 21481 18914 21516 18978
rect 21371 18897 21516 18914
rect 26221 18975 26417 18991
rect 26221 18903 26281 18975
rect 26370 18903 26417 18975
rect 26221 18887 26417 18903
rect 31024 18969 31249 18988
rect 31024 18911 31080 18969
rect 31192 18911 31249 18969
rect 31024 18894 31249 18911
rect 37099 18978 37284 18996
rect 37099 18909 37151 18978
rect 37227 18909 37284 18978
rect 37099 18894 37284 18909
rect 3807 18136 4033 18157
rect 336 18072 560 18097
rect 336 18005 392 18072
rect 505 18005 560 18072
rect 3807 18059 3863 18136
rect 3977 18059 4033 18136
rect 3807 18031 4033 18059
rect 8625 18139 8848 18176
rect 8625 18055 8680 18139
rect 8792 18055 8848 18139
rect 8625 18028 8848 18055
rect 13840 18138 14050 18175
rect 13840 18070 13888 18138
rect 14002 18070 14050 18138
rect 13840 18039 14050 18070
rect 18228 18144 18387 18174
rect 18228 18065 18269 18144
rect 18349 18065 18387 18144
rect 18228 18041 18387 18065
rect 23408 18143 23632 18167
rect 23408 18068 23464 18143
rect 23575 18068 23632 18143
rect 23408 18032 23632 18068
rect 27833 18139 28057 18167
rect 27833 18066 27889 18139
rect 28002 18066 28057 18139
rect 27833 18031 28057 18066
rect 32985 18117 33201 18139
rect 32985 18053 33038 18117
rect 33154 18053 33201 18117
rect 32985 18031 33201 18053
rect 35758 18127 35923 18147
rect 35758 18068 35784 18127
rect 35896 18068 35923 18127
rect 35758 18043 35923 18068
rect 336 17979 560 18005
rect 441 17675 524 17685
rect 212 17616 301 17621
rect 212 17561 231 17616
rect 284 17561 301 17616
rect 441 17618 451 17675
rect 514 17618 524 17675
rect 441 17608 524 17618
rect 212 17555 301 17561
rect 212 17545 294 17555
rect -1344 17489 294 17545
rect -1344 15921 -1007 17489
rect 2128 17300 2352 17315
rect 2128 17214 2184 17300
rect 2296 17214 2352 17300
rect 2128 17195 2352 17214
rect 6830 17291 7055 17313
rect 6830 17221 6888 17291
rect 7000 17221 7055 17291
rect 6830 17195 7055 17221
rect 11704 17282 11928 17314
rect 11704 17212 11761 17282
rect 11872 17212 11928 17282
rect 11704 17195 11928 17212
rect 16564 17278 16708 17295
rect 16564 17219 16599 17278
rect 16671 17219 16708 17278
rect 16564 17199 16708 17219
rect 21380 17285 21525 17299
rect 21380 17212 21407 17285
rect 21487 17212 21525 17285
rect 21380 17201 21525 17212
rect 26223 17285 26419 17304
rect 26223 17214 26270 17285
rect 26369 17214 26419 17285
rect 26223 17200 26419 17214
rect 31024 17279 31248 17294
rect 31024 17221 31080 17279
rect 31192 17221 31248 17279
rect 31024 17204 31248 17221
rect 37099 17289 37264 17304
rect 37099 17220 37143 17289
rect 37219 17220 37264 17289
rect 37099 17208 37264 17220
rect 2128 16181 2352 16203
rect 2128 16117 2184 16181
rect 2296 16117 2352 16181
rect 2128 16083 2352 16117
rect 6832 16173 7057 16200
rect 6832 16104 6887 16173
rect 7000 16104 7057 16173
rect 6832 16082 7057 16104
rect 11704 16180 11929 16203
rect 11704 16110 11762 16180
rect 11873 16110 11929 16180
rect 11704 16083 11929 16110
rect 16560 16175 16704 16193
rect 16560 16114 16588 16175
rect 16667 16114 16704 16175
rect 16560 16097 16704 16114
rect 21366 16181 21537 16197
rect 21366 16108 21411 16181
rect 21491 16108 21537 16181
rect 21366 16093 21537 16108
rect 26234 16176 26408 16192
rect 26234 16105 26271 16176
rect 26370 16105 26408 16176
rect 26234 16088 26408 16105
rect 31024 16171 31248 16187
rect 31024 16115 31080 16171
rect 31192 16115 31248 16171
rect 31024 16097 31248 16115
rect 37096 16175 37261 16191
rect 37096 16111 37144 16175
rect 37218 16111 37261 16175
rect 37096 16095 37261 16111
rect -1344 15849 512 15921
rect -1344 12051 -1007 15849
rect 440 15793 512 15849
rect 432 15779 519 15793
rect 432 15724 450 15779
rect 505 15724 519 15779
rect 432 15710 519 15724
rect 335 15321 561 15359
rect 335 15254 378 15321
rect 513 15254 561 15321
rect 335 15232 561 15254
rect 3808 15332 4034 15373
rect 3808 15255 3863 15332
rect 3977 15255 4034 15332
rect 3808 15231 4034 15255
rect 8624 15343 8849 15372
rect 8624 15249 8679 15343
rect 8791 15249 8849 15343
rect 8624 15218 8849 15249
rect 13846 15338 14056 15369
rect 13846 15263 13887 15338
rect 14008 15263 14056 15338
rect 13846 15233 14056 15263
rect 18235 15336 18394 15369
rect 18235 15261 18267 15336
rect 18351 15261 18394 15336
rect 18235 15236 18394 15261
rect 23409 15324 23633 15368
rect 23409 15258 23462 15324
rect 23577 15258 23633 15324
rect 23409 15233 23633 15258
rect 27832 15334 28056 15371
rect 27832 15263 27888 15334
rect 28000 15263 28056 15334
rect 27832 15235 28056 15263
rect 32988 15339 33204 15360
rect 32988 15269 33040 15339
rect 33152 15269 33204 15339
rect 32988 15252 33204 15269
rect 35755 15333 35920 15357
rect 35755 15274 35784 15333
rect 35896 15274 35920 15333
rect 35755 15253 35920 15274
rect 2128 14495 2352 14515
rect 2128 14425 2184 14495
rect 2296 14425 2352 14495
rect 2128 14395 2352 14425
rect 6832 14489 7056 14515
rect 6832 14420 6888 14489
rect 7001 14420 7056 14489
rect 6832 14395 7056 14420
rect 11704 14494 11929 14515
rect 11704 14418 11760 14494
rect 11873 14418 11929 14494
rect 11704 14395 11929 14418
rect 16555 14478 16714 14499
rect 16555 14417 16592 14478
rect 16671 14417 16714 14478
rect 16555 14401 16714 14417
rect 21358 14481 21529 14504
rect 21358 14410 21397 14481
rect 21484 14410 21529 14481
rect 21358 14400 21529 14410
rect 26228 14483 26402 14503
rect 26228 14414 26265 14483
rect 26371 14414 26402 14483
rect 26228 14399 26402 14414
rect 31024 14479 31249 14498
rect 31024 14423 31080 14479
rect 31192 14423 31249 14479
rect 31024 14406 31249 14423
rect 37105 14489 37272 14508
rect 37105 14425 37150 14489
rect 37224 14425 37272 14489
rect 37105 14405 37272 14425
rect 2128 13383 2352 13403
rect 2128 13310 2184 13383
rect 2296 13310 2352 13383
rect 2128 13283 2352 13310
rect 6832 13374 7056 13403
rect 6832 13305 6885 13374
rect 7001 13305 7056 13374
rect 6832 13283 7056 13305
rect 11704 13384 11929 13402
rect 11704 13308 11760 13384
rect 11873 13308 11929 13384
rect 11704 13283 11929 13308
rect 16547 13372 16706 13392
rect 16547 13308 16594 13372
rect 16668 13308 16706 13372
rect 16547 13294 16706 13308
rect 21375 13376 21526 13393
rect 21375 13305 21406 13376
rect 21493 13305 21526 13376
rect 21375 13288 21526 13305
rect 26228 13380 26410 13396
rect 26228 13311 26267 13380
rect 26373 13311 26410 13380
rect 26228 13292 26410 13311
rect 31024 13370 31249 13390
rect 31024 13310 31080 13370
rect 31192 13310 31249 13370
rect 31024 13298 31249 13310
rect 37107 13376 37274 13394
rect 37107 13308 37148 13376
rect 37226 13308 37274 13376
rect 37107 13291 37274 13308
rect 3807 12535 4033 12574
rect 363 12463 532 12498
rect 363 12402 396 12463
rect 501 12402 532 12463
rect 3807 12464 3864 12535
rect 3977 12464 4033 12535
rect 3807 12432 4033 12464
rect 8624 12549 8849 12574
rect 8624 12455 8681 12549
rect 8793 12455 8849 12549
rect 8624 12429 8849 12455
rect 13830 12535 14058 12579
rect 13830 12460 13885 12535
rect 14006 12460 14058 12535
rect 13830 12432 14058 12460
rect 18216 12530 18394 12566
rect 18216 12455 18268 12530
rect 18352 12455 18394 12530
rect 18216 12431 18394 12455
rect 23408 12526 23633 12555
rect 23408 12460 23462 12526
rect 23577 12460 23633 12526
rect 23408 12432 23633 12460
rect 27833 12527 28055 12559
rect 27833 12456 27889 12527
rect 28001 12456 28055 12527
rect 27833 12431 28055 12456
rect 33004 12535 33183 12558
rect 33004 12465 33040 12535
rect 33152 12465 33183 12535
rect 33004 12445 33183 12465
rect 35750 12524 35932 12542
rect 35750 12465 35784 12524
rect 35896 12465 35932 12524
rect 35750 12442 35932 12465
rect 363 12379 532 12402
rect 428 12051 523 12054
rect -1344 12043 523 12051
rect -1344 11987 450 12043
rect 507 11987 523 12043
rect -1344 11983 523 11987
rect -1344 10098 -1007 11983
rect 428 11975 523 11983
rect 2128 11700 2352 11715
rect 2128 11616 2184 11700
rect 2296 11616 2352 11700
rect 2128 11595 2352 11616
rect 6832 11684 7056 11714
rect 6832 11615 6886 11684
rect 7002 11615 7056 11684
rect 6832 11594 7056 11615
rect 11704 11686 11929 11714
rect 11704 11611 11760 11686
rect 11872 11611 11929 11686
rect 11704 11595 11929 11611
rect 16567 11681 16716 11697
rect 16567 11617 16601 11681
rect 16675 11617 16716 11681
rect 16567 11603 16716 11617
rect 21365 11686 21516 11704
rect 21365 11610 21397 11686
rect 21483 11610 21516 11686
rect 21365 11599 21516 11610
rect 26230 11687 26412 11703
rect 26230 11611 26278 11687
rect 26367 11611 26412 11687
rect 26230 11599 26412 11611
rect 31024 11685 31248 11698
rect 31024 11625 31080 11685
rect 31192 11625 31248 11685
rect 31024 11610 31248 11625
rect 37094 11686 37270 11704
rect 37094 11618 37146 11686
rect 37224 11618 37270 11686
rect 37094 11603 37270 11618
rect 31025 10736 31249 10824
rect 2128 10581 2352 10603
rect 2128 10503 2184 10581
rect 2296 10503 2352 10581
rect 2128 10483 2352 10503
rect 6831 10576 7055 10602
rect 6831 10505 6887 10576
rect 7001 10505 7055 10576
rect 6831 10482 7055 10505
rect 11704 10583 11928 10603
rect 11704 10508 11760 10583
rect 11872 10508 11928 10583
rect 11704 10483 11928 10508
rect 16560 10574 16709 10592
rect 16560 10512 16593 10574
rect 16669 10512 16709 10574
rect 16560 10498 16709 10512
rect 21357 10576 21525 10591
rect 21357 10500 21402 10576
rect 21488 10500 21525 10576
rect 21357 10489 21525 10500
rect 26228 10582 26415 10596
rect 26228 10506 26277 10582
rect 26366 10506 26415 10582
rect 26228 10489 26415 10506
rect 31024 10574 31248 10590
rect 31024 10518 31080 10574
rect 31193 10518 31248 10574
rect 31024 10502 31248 10518
rect 37093 10579 37269 10594
rect 37093 10506 37137 10579
rect 37219 10506 37269 10579
rect 37093 10493 37269 10506
rect 447 10178 530 10188
rect 447 10123 461 10178
rect 516 10123 530 10178
rect 447 10115 530 10123
rect 447 10098 524 10115
rect -1344 10026 524 10098
rect -1344 6478 -1007 10026
rect 452 10025 524 10026
rect 336 9719 503 9744
rect 336 9654 368 9719
rect 474 9654 503 9719
rect 336 9632 503 9654
rect 3808 9741 4034 9767
rect 3808 9670 3863 9741
rect 3976 9670 4034 9741
rect 3808 9632 4034 9670
rect 8622 9730 8847 9762
rect 8622 9647 8680 9730
rect 8794 9647 8847 9730
rect 8622 9617 8847 9647
rect 13830 9735 14058 9780
rect 13830 9663 13887 9735
rect 14004 9663 14058 9735
rect 13830 9633 14058 9663
rect 18213 9735 18391 9766
rect 18213 9655 18265 9735
rect 18353 9655 18391 9735
rect 18213 9631 18391 9655
rect 23407 9726 23632 9763
rect 23407 9663 23463 9726
rect 23578 9663 23632 9726
rect 23407 9640 23632 9663
rect 27833 9733 28055 9762
rect 27833 9663 27888 9733
rect 28000 9663 28055 9733
rect 27833 9634 28055 9663
rect 33003 9732 33182 9760
rect 33003 9666 33031 9732
rect 33143 9666 33182 9732
rect 33003 9647 33182 9666
rect 35745 9732 35927 9755
rect 35745 9674 35784 9732
rect 35896 9674 35927 9732
rect 35745 9655 35927 9674
rect 334 9278 419 9288
rect 334 9214 344 9278
rect 408 9214 419 9278
rect 334 9203 419 9214
rect 2128 8893 2352 8915
rect 2128 8813 2184 8893
rect 2296 8813 2352 8893
rect 2128 8795 2352 8813
rect 6833 8885 7057 8913
rect 6833 8814 6886 8885
rect 7000 8814 7057 8885
rect 6833 8795 7057 8814
rect 11704 8889 11928 8914
rect 11704 8811 11760 8889
rect 11872 8811 11928 8889
rect 11704 8794 11928 8811
rect 16551 8878 16727 8900
rect 16551 8816 16598 8878
rect 16674 8816 16727 8878
rect 16551 8802 16727 8816
rect 21357 8885 21525 8904
rect 21357 8811 21397 8885
rect 21484 8811 21525 8885
rect 21357 8802 21525 8811
rect 26223 8886 26410 8907
rect 26223 8811 26265 8886
rect 26364 8811 26410 8886
rect 26223 8800 26410 8811
rect 31033 8882 31231 8900
rect 31033 8826 31079 8882
rect 31192 8826 31231 8882
rect 31033 8807 31231 8826
rect 37092 8885 37270 8901
rect 37092 8812 37142 8885
rect 37224 8812 37270 8885
rect 37092 8802 37270 8812
rect 2128 7784 2352 7803
rect 2128 7714 2184 7784
rect 2296 7714 2352 7784
rect 2128 7683 2352 7714
rect 6832 7773 7056 7802
rect 6832 7708 6888 7773
rect 7000 7708 7056 7773
rect 6832 7684 7056 7708
rect 11704 7781 11928 7802
rect 11704 7703 11760 7781
rect 11872 7703 11928 7781
rect 11704 7683 11928 7703
rect 16540 7772 16716 7791
rect 16540 7706 16589 7772
rect 16670 7706 16716 7772
rect 16540 7693 16716 7706
rect 21363 7779 21532 7793
rect 21363 7705 21404 7779
rect 21491 7705 21532 7779
rect 21363 7689 21532 7705
rect 26231 7783 26414 7796
rect 26231 7708 26273 7783
rect 26372 7708 26414 7783
rect 26231 7693 26414 7708
rect 31031 7772 31229 7790
rect 31031 7716 31079 7772
rect 31192 7716 31229 7772
rect 31031 7697 31229 7716
rect 37097 7779 37275 7794
rect 37097 7711 37144 7779
rect 37228 7711 37275 7779
rect 37097 7695 37275 7711
rect 3807 6935 4033 6967
rect 337 6874 561 6900
rect 337 6805 390 6874
rect 505 6805 561 6874
rect 3807 6854 3863 6935
rect 3977 6854 4033 6935
rect 3807 6832 4033 6854
rect 8623 6928 8848 6965
rect 8623 6849 8679 6928
rect 8791 6849 8848 6928
rect 8623 6824 8848 6849
rect 13832 6938 14058 6973
rect 13832 6866 13886 6938
rect 14003 6866 14058 6938
rect 13832 6838 14058 6866
rect 18225 6956 18392 6977
rect 18225 6876 18263 6956
rect 18351 6876 18392 6956
rect 18225 6855 18392 6876
rect 23406 6928 23634 6962
rect 23406 6865 23462 6928
rect 23577 6865 23634 6928
rect 23406 6834 23634 6865
rect 27831 6939 28053 6967
rect 27831 6869 27887 6939
rect 27999 6869 28053 6939
rect 27831 6832 28053 6869
rect 33009 6930 33190 6951
rect 33009 6864 33041 6930
rect 33153 6864 33190 6930
rect 33009 6842 33190 6864
rect 35737 6921 35937 6945
rect 35737 6863 35784 6921
rect 35896 6863 35937 6921
rect 35737 6839 35937 6863
rect 337 6779 561 6805
rect 320 6478 406 6482
rect -1344 6473 406 6478
rect -1344 6421 334 6473
rect 389 6421 406 6473
rect -1344 6415 406 6421
rect -1344 4735 -1007 6415
rect 320 6408 406 6415
rect 544 6479 628 6489
rect 544 6416 554 6479
rect 618 6416 628 6479
rect 544 6406 628 6416
rect 2128 6088 2352 6115
rect 2128 6012 2184 6088
rect 2296 6012 2352 6088
rect 2128 5995 2352 6012
rect 6832 6081 7056 6115
rect 6832 6016 6888 6081
rect 7000 6016 7056 6081
rect 6832 5995 7056 6016
rect 11703 6089 11927 6114
rect 11703 6016 11761 6089
rect 11874 6016 11927 6089
rect 11703 5995 11927 6016
rect 16558 6082 16730 6104
rect 16558 6016 16593 6082
rect 16674 6016 16730 6082
rect 16558 5998 16730 6016
rect 21359 6083 21528 6105
rect 21359 6011 21400 6083
rect 21485 6011 21528 6083
rect 21359 6001 21528 6011
rect 26232 6090 26415 6102
rect 26232 6010 26275 6090
rect 26367 6010 26415 6090
rect 26232 5999 26415 6010
rect 31049 6082 31220 6098
rect 31049 6026 31080 6082
rect 31193 6026 31220 6082
rect 31049 6009 31220 6026
rect 37090 6083 37270 6101
rect 37090 6015 37140 6083
rect 37224 6015 37270 6083
rect 37090 6002 37270 6015
rect 2128 4984 2353 5003
rect 2128 4910 2184 4984
rect 2296 4910 2353 4984
rect 2128 4883 2353 4910
rect 6832 4974 7056 5003
rect 6832 4903 6888 4974
rect 7001 4903 7056 4974
rect 6832 4883 7056 4903
rect 11704 4980 11929 5002
rect 11704 4907 11759 4980
rect 11872 4907 11929 4980
rect 11704 4883 11929 4907
rect 16545 4976 16717 4993
rect 16545 4906 16589 4976
rect 16672 4906 16717 4976
rect 16545 4887 16717 4906
rect 21375 4974 21532 4993
rect 21375 4902 21408 4974
rect 21493 4902 21532 4974
rect 21375 4887 21532 4902
rect 26242 4980 26415 4996
rect 26242 4900 26281 4980
rect 26373 4900 26415 4980
rect 31050 4977 31221 4990
rect 31050 4921 31080 4977
rect 31192 4921 31221 4977
rect 31050 4901 31221 4921
rect 37100 4976 37280 4992
rect 37100 4910 37140 4976
rect 37228 4910 37280 4976
rect 26242 4886 26415 4900
rect 37100 4893 37280 4910
rect -1344 4663 618 4735
rect -1344 2800 -1007 4663
rect 546 4590 618 4663
rect 536 4577 626 4590
rect 536 4523 557 4577
rect 611 4523 626 4577
rect 536 4506 626 4523
rect 336 4141 561 4200
rect 336 4062 390 4141
rect 507 4062 561 4141
rect 336 4028 561 4062
rect 3808 4139 4032 4172
rect 3808 4058 3863 4139
rect 3977 4058 4032 4139
rect 3808 4031 4032 4058
rect 8624 4129 8849 4164
rect 8624 4052 8680 4129
rect 8793 4052 8849 4129
rect 8624 4025 8849 4052
rect 13831 4135 14057 4166
rect 13831 4060 13887 4135
rect 14000 4060 14057 4135
rect 13831 4033 14057 4060
rect 18222 4141 18389 4170
rect 18222 4066 18267 4141
rect 18360 4066 18389 4141
rect 18222 4048 18389 4066
rect 23407 4127 23635 4161
rect 23407 4056 23460 4127
rect 23576 4056 23635 4127
rect 23407 4033 23635 4056
rect 27834 4123 28056 4160
rect 27834 4050 27887 4123
rect 28001 4050 28056 4123
rect 27834 4025 28056 4050
rect 32997 4136 33178 4158
rect 32997 4072 33030 4136
rect 33139 4072 33178 4136
rect 32997 4049 33178 4072
rect 35742 4130 35942 4159
rect 35742 4074 35783 4130
rect 35896 4074 35942 4130
rect 35742 4053 35942 4074
rect 318 3677 401 3687
rect 318 3617 328 3677
rect 391 3617 401 3677
rect 318 3607 401 3617
rect 2128 3293 2352 3315
rect 2128 3214 2184 3293
rect 2296 3214 2352 3293
rect 2128 3195 2352 3214
rect 6832 3288 7056 3314
rect 6832 3217 6888 3288
rect 7001 3217 7056 3288
rect 6832 3194 7056 3217
rect 11701 3284 11926 3314
rect 11701 3209 11757 3284
rect 11875 3209 11926 3284
rect 11701 3195 11926 3209
rect 16560 3288 16719 3302
rect 16560 3218 16594 3288
rect 16677 3218 16719 3288
rect 16560 3202 16719 3218
rect 21371 3283 21528 3303
rect 21371 3212 21401 3283
rect 21486 3212 21528 3283
rect 21371 3197 21528 3212
rect 26229 3290 26402 3309
rect 26229 3210 26264 3290
rect 26360 3210 26402 3290
rect 26229 3199 26402 3210
rect 31051 3278 31233 3299
rect 31051 3222 31080 3278
rect 31192 3222 31233 3278
rect 31051 3204 31233 3222
rect 37093 3285 37278 3305
rect 37093 3219 37137 3285
rect 37225 3219 37278 3285
rect 37093 3206 37278 3219
rect 2128 2172 2352 2203
rect 2128 2104 2184 2172
rect 2296 2104 2352 2172
rect 2128 2083 2352 2104
rect 6832 2173 7056 2204
rect 6832 2104 6887 2173
rect 7001 2104 7056 2173
rect 6832 2084 7056 2104
rect 11702 2181 11929 2200
rect 11702 2106 11758 2181
rect 11876 2106 11929 2181
rect 11702 2085 11929 2106
rect 16553 2177 16712 2194
rect 16553 2104 16595 2177
rect 16675 2104 16712 2177
rect 16553 2094 16712 2104
rect 21376 2174 21524 2196
rect 21376 2103 21403 2174
rect 21488 2103 21524 2174
rect 21376 2084 21524 2103
rect 26227 2179 26412 2195
rect 26227 2099 26276 2179
rect 26372 2099 26412 2179
rect 31046 2178 31228 2194
rect 31046 2117 31079 2178
rect 31193 2117 31228 2178
rect 31046 2099 31228 2117
rect 26227 2088 26412 2099
rect 3808 1332 4032 1378
rect 3808 1265 3864 1332
rect 3976 1265 4032 1332
rect 3808 1232 4032 1265
rect 8625 1334 8849 1364
rect 8625 1257 8679 1334
rect 8792 1257 8849 1334
rect 8625 1231 8849 1257
rect 13834 1328 14055 1363
rect 13834 1255 13872 1328
rect 14002 1255 14055 1328
rect 13834 1219 14055 1255
rect 18198 1335 18424 1361
rect 18198 1260 18262 1335
rect 18355 1260 18424 1335
rect 18198 1233 18424 1260
rect 23409 1342 23632 1368
rect 23409 1271 23462 1342
rect 23578 1271 23632 1342
rect 23409 1233 23632 1271
rect 27832 1330 28059 1357
rect 27832 1257 27887 1330
rect 28001 1257 28059 1330
rect 27832 1233 28059 1257
rect 33008 1329 33186 1356
rect 33008 1265 33043 1329
rect 33152 1265 33186 1329
rect 33008 1241 33186 1265
rect 2128 489 2352 515
rect 2128 416 2184 489
rect 2296 416 2352 489
rect 2128 395 2352 416
rect 6831 487 7057 515
rect 6831 418 6887 487
rect 7001 418 7057 487
rect 6831 395 7057 418
rect 11704 487 11931 511
rect 11704 410 11760 487
rect 11872 410 11931 487
rect 11704 396 11931 410
rect 16529 485 16723 502
rect 16529 412 16588 485
rect 16668 412 16723 485
rect 16529 401 16723 412
rect 21369 480 21517 507
rect 21369 408 21402 480
rect 21481 408 21517 480
rect 21369 395 21517 408
rect 26229 483 26414 505
rect 26229 406 26275 483
rect 26363 406 26414 483
rect 26229 398 26414 406
rect 31041 482 31228 504
rect 31041 421 31079 482
rect 31193 421 31228 482
rect 31041 402 31228 421
<< via2 >>
rect 472 24324 530 24380
rect 391 22657 504 22733
rect 3881 22614 3971 22672
rect 8680 23169 8793 23243
rect 13888 23184 13944 23240
rect 10358 22848 10418 22850
rect 10358 22794 10361 22848
rect 10361 22794 10415 22848
rect 10415 22794 10418 22848
rect 10358 22792 10418 22794
rect 18283 23184 18339 23240
rect 23493 23184 23549 23240
rect 27862 23179 28000 23251
rect 35783 26137 35896 26199
rect 37139 25335 37230 25411
rect 35784 25176 35897 25238
rect 37137 24378 37228 24454
rect 35784 24221 35896 24283
rect 37140 23426 37220 23495
rect 29788 22792 29852 22852
rect 35784 23238 35896 23300
rect 11761 22389 11874 22465
rect 16605 22400 16661 22456
rect 21421 22400 21477 22456
rect 26292 22400 26348 22456
rect 31111 22400 31167 22456
rect 37137 22449 37216 22518
rect 3862 22224 3923 22226
rect 3862 22172 3865 22224
rect 3865 22172 3920 22224
rect 3920 22172 3923 22224
rect 3862 22170 3923 22172
rect 2184 21703 2296 21777
rect 6887 21698 7001 21776
rect 11760 21700 11873 21782
rect 16593 21710 16683 21769
rect 21412 21709 21490 21773
rect 26264 21706 26375 21776
rect 31080 21714 31193 21771
rect 37146 21707 37224 21773
rect 467 21377 528 21380
rect 467 21325 470 21377
rect 470 21325 525 21377
rect 525 21325 528 21377
rect 467 21323 528 21325
rect 392 20849 505 20925
rect 3864 20871 3976 20940
rect 8678 20855 8793 20940
rect 13889 20866 14003 20934
rect 18268 20864 18348 20943
rect 23462 20862 23576 20944
rect 27887 20864 28000 20937
rect 33039 20874 33155 20938
rect 35784 20869 35896 20928
rect 2184 20019 2296 20085
rect 6888 20014 7000 20091
rect 11760 20016 11872 20098
rect 16583 20022 16673 20081
rect 21409 20021 21486 20085
rect 26277 20017 26366 20089
rect 31079 20020 31192 20077
rect 37145 20023 37223 20089
rect 2184 18907 2296 18973
rect 6888 18901 7000 18976
rect 11760 18904 11872 18986
rect 16593 18910 16665 18969
rect 21404 18914 21481 18978
rect 26281 18903 26370 18975
rect 31080 18911 31192 18969
rect 37151 18909 37227 18978
rect 392 18005 505 18072
rect 3863 18059 3977 18136
rect 8680 18055 8792 18139
rect 13888 18070 14002 18138
rect 18269 18065 18349 18144
rect 23464 18068 23575 18143
rect 27889 18066 28002 18139
rect 33038 18053 33154 18117
rect 35784 18068 35896 18127
rect 451 17673 514 17675
rect 451 17621 454 17673
rect 454 17621 510 17673
rect 510 17621 514 17673
rect 451 17618 514 17621
rect 2184 17214 2296 17300
rect 6888 17221 7000 17291
rect 11761 17212 11872 17282
rect 16599 17219 16671 17278
rect 21407 17212 21487 17285
rect 26270 17214 26369 17285
rect 31080 17221 31192 17279
rect 37143 17220 37219 17289
rect 2184 16117 2296 16181
rect 6887 16104 7000 16173
rect 11762 16110 11873 16180
rect 16588 16114 16667 16175
rect 21411 16108 21491 16181
rect 26271 16105 26370 16176
rect 31080 16115 31192 16171
rect 37144 16111 37218 16175
rect 378 15254 513 15321
rect 3863 15255 3977 15332
rect 8679 15249 8791 15343
rect 13887 15263 14008 15338
rect 18267 15261 18351 15336
rect 23462 15258 23577 15324
rect 27888 15263 28000 15334
rect 33040 15269 33152 15339
rect 35784 15274 35896 15333
rect 2184 14425 2296 14495
rect 6888 14420 7001 14489
rect 11760 14418 11873 14494
rect 16592 14417 16671 14478
rect 21397 14410 21484 14481
rect 26265 14414 26371 14483
rect 31080 14423 31192 14479
rect 37150 14425 37224 14489
rect 2184 13310 2296 13383
rect 6885 13305 7001 13374
rect 11760 13308 11873 13384
rect 16594 13308 16668 13372
rect 21406 13305 21493 13376
rect 26267 13311 26373 13380
rect 31080 13310 31192 13370
rect 37148 13308 37226 13376
rect 396 12402 501 12463
rect 3864 12464 3977 12535
rect 8681 12455 8793 12549
rect 13885 12460 14006 12535
rect 18268 12455 18352 12530
rect 23462 12460 23577 12526
rect 27889 12456 28001 12527
rect 33040 12465 33152 12535
rect 35784 12465 35896 12524
rect 2184 11616 2296 11700
rect 6886 11615 7002 11684
rect 11760 11611 11872 11686
rect 16601 11617 16675 11681
rect 21397 11610 21483 11686
rect 26278 11611 26367 11687
rect 31080 11625 31192 11685
rect 37146 11618 37224 11686
rect 2184 10503 2296 10581
rect 6887 10505 7001 10576
rect 11760 10508 11872 10583
rect 16593 10512 16669 10574
rect 21402 10500 21488 10576
rect 26277 10506 26366 10582
rect 31080 10573 31193 10574
rect 31080 10518 31193 10573
rect 37137 10506 37219 10579
rect 368 9654 474 9719
rect 3863 9670 3976 9741
rect 8680 9647 8794 9730
rect 13887 9663 14004 9735
rect 18265 9655 18353 9735
rect 23463 9663 23578 9726
rect 27888 9663 28000 9733
rect 33031 9666 33143 9732
rect 35784 9674 35896 9732
rect 344 9274 408 9278
rect 344 9217 347 9274
rect 347 9217 404 9274
rect 404 9217 408 9274
rect 344 9214 408 9217
rect 2184 8813 2296 8893
rect 6886 8814 7000 8885
rect 11760 8811 11872 8889
rect 16598 8816 16674 8878
rect 21397 8811 21484 8885
rect 26265 8811 26364 8886
rect 31079 8826 31192 8882
rect 37142 8812 37224 8885
rect 2184 7714 2296 7784
rect 6888 7708 7000 7773
rect 11760 7703 11872 7781
rect 16589 7706 16670 7772
rect 21404 7705 21491 7779
rect 26273 7708 26372 7783
rect 31079 7716 31192 7772
rect 37144 7711 37228 7779
rect 390 6805 505 6874
rect 3863 6854 3977 6935
rect 8679 6849 8791 6928
rect 13886 6866 14003 6938
rect 18263 6876 18351 6956
rect 23462 6865 23577 6928
rect 27887 6869 27999 6939
rect 33041 6864 33153 6930
rect 35784 6863 35896 6921
rect 554 6416 618 6479
rect 2184 6012 2296 6088
rect 6888 6016 7000 6081
rect 11761 6016 11874 6089
rect 16593 6016 16674 6082
rect 21400 6011 21485 6083
rect 26275 6010 26367 6090
rect 31080 6026 31193 6082
rect 37140 6015 37224 6083
rect 2184 4910 2296 4984
rect 6888 4903 7001 4974
rect 11759 4907 11872 4980
rect 16589 4906 16672 4976
rect 21408 4902 21493 4974
rect 26281 4900 26373 4980
rect 31080 4921 31192 4977
rect 37140 4910 37228 4976
rect 390 4062 507 4141
rect 3863 4058 3977 4139
rect 8680 4052 8793 4129
rect 13887 4060 14000 4135
rect 18267 4066 18360 4141
rect 23460 4056 23576 4127
rect 27887 4050 28001 4123
rect 33030 4072 33139 4136
rect 35783 4074 35896 4130
rect 328 3674 391 3677
rect 328 3620 333 3674
rect 333 3620 388 3674
rect 388 3620 391 3674
rect 328 3617 391 3620
rect 2184 3214 2296 3293
rect 6888 3217 7001 3288
rect 11757 3209 11875 3284
rect 16594 3218 16677 3288
rect 21401 3212 21486 3283
rect 26264 3210 26360 3290
rect 31080 3222 31192 3278
rect 37137 3219 37225 3285
rect 2184 2104 2296 2172
rect 6887 2104 7001 2173
rect 11758 2106 11876 2181
rect 16595 2104 16675 2177
rect 21403 2103 21488 2174
rect 26276 2099 26372 2179
rect 31079 2117 31193 2178
rect 3864 1265 3976 1332
rect 8679 1257 8792 1334
rect 13872 1255 14002 1328
rect 18262 1260 18355 1335
rect 23462 1271 23578 1342
rect 27887 1257 28001 1330
rect 33043 1265 33152 1329
rect 2184 416 2296 489
rect 6887 418 7001 487
rect 11760 410 11872 487
rect 16588 412 16668 485
rect 21402 408 21481 480
rect 26275 406 26363 483
rect 31079 421 31193 482
<< metal3 >>
rect 40053 36415 40873 37242
rect 3163 35114 3983 35941
rect 3416 30816 3754 35114
rect 16944 35100 17764 35927
rect 3414 30408 3754 30816
rect 3414 26824 3752 30408
rect -1736 26600 3752 26824
rect -1736 25396 -1400 26600
rect 3414 26543 3752 26600
rect 17191 26880 17527 35100
rect 40264 35078 40597 36415
rect 17191 26544 17528 26880
rect 40264 26712 40599 35078
rect 17191 26543 17527 26544
rect -1736 21384 -1399 25396
rect 6473 24585 7469 24588
rect 17248 24585 17472 26543
rect 40264 26376 40600 26712
rect 35728 26199 35952 26214
rect 35728 26137 35783 26199
rect 35896 26137 35952 26199
rect 35728 26113 35952 26137
rect 37095 25411 37276 25429
rect 37095 25335 37139 25411
rect 37230 25335 37276 25411
rect 37095 25320 37276 25335
rect 35750 25238 35928 25254
rect 35750 25176 35784 25238
rect 35897 25176 35928 25238
rect 35750 25154 35928 25176
rect 224 24380 30464 24585
rect 224 24324 472 24380
rect 530 24324 30464 24380
rect 37085 24454 37283 24467
rect 37085 24378 37137 24454
rect 37228 24378 37283 24454
rect 37085 24368 37283 24378
rect 224 24248 30464 24324
rect 35748 24283 35926 24295
rect 2022 24247 2541 24248
rect 336 22733 562 22762
rect 336 22657 391 22733
rect 504 22657 562 22733
rect 336 22628 562 22657
rect 3633 22237 3710 24248
rect 8624 23243 8847 23275
rect 8624 23169 8680 23243
rect 8793 23169 8847 23243
rect 8624 23154 8847 23169
rect 10352 22860 10424 24248
rect 11310 24247 12106 24248
rect 16409 24247 16979 24248
rect 27843 23251 28014 23274
rect 13878 23240 13954 23250
rect 13878 23184 13888 23240
rect 13944 23184 13954 23240
rect 13878 23174 13954 23184
rect 18273 23240 18349 23250
rect 18273 23184 18283 23240
rect 18339 23184 18349 23240
rect 18273 23174 18349 23184
rect 23483 23240 23559 23250
rect 23483 23184 23493 23240
rect 23549 23184 23559 23240
rect 23483 23174 23559 23184
rect 27843 23179 27862 23251
rect 28000 23179 28014 23251
rect 27843 23158 28014 23179
rect 29782 22862 29854 24248
rect 35748 24221 35784 24283
rect 35896 24221 35926 24283
rect 35748 24195 35926 24221
rect 37085 23495 37283 23510
rect 37085 23426 37140 23495
rect 37220 23426 37283 23495
rect 37085 23411 37283 23426
rect 35739 23300 35940 23321
rect 35739 23238 35784 23300
rect 35896 23238 35940 23300
rect 35739 23218 35940 23238
rect 10348 22850 10428 22860
rect 10348 22792 10358 22850
rect 10418 22792 10428 22850
rect 10348 22782 10428 22792
rect 29778 22852 29862 22862
rect 29778 22792 29788 22852
rect 29852 22792 29862 22852
rect 29778 22782 29862 22792
rect 3836 22672 4021 22707
rect 3836 22614 3881 22672
rect 3971 22614 4021 22672
rect 3836 22586 4021 22614
rect 37101 22518 37264 22537
rect 11727 22465 11904 22491
rect 11727 22389 11761 22465
rect 11874 22389 11904 22465
rect 16595 22456 16671 22466
rect 16595 22400 16605 22456
rect 16661 22400 16671 22456
rect 16595 22390 16671 22400
rect 21411 22456 21487 22466
rect 21411 22400 21421 22456
rect 21477 22400 21487 22456
rect 21411 22390 21487 22400
rect 26282 22456 26358 22466
rect 26282 22400 26292 22456
rect 26348 22400 26358 22456
rect 26282 22390 26358 22400
rect 31101 22456 31177 22466
rect 31101 22400 31111 22456
rect 31167 22400 31177 22456
rect 37101 22449 37137 22518
rect 37217 22449 37264 22518
rect 37101 22436 37264 22449
rect 31101 22390 31177 22400
rect 11727 22369 11904 22389
rect 3633 22226 3934 22237
rect 3633 22170 3862 22226
rect 3923 22170 3934 22226
rect 3633 22160 3934 22170
rect 3851 22159 3934 22160
rect 2128 21777 2352 21803
rect 2128 21703 2184 21777
rect 2296 21703 2352 21777
rect 2128 21683 2352 21703
rect 6832 21776 7056 21803
rect 6832 21698 6887 21776
rect 7001 21698 7056 21776
rect 6832 21683 7056 21698
rect 11704 21782 11928 21803
rect 11704 21700 11760 21782
rect 11873 21700 11928 21782
rect 11704 21683 11928 21700
rect 16520 21769 16744 21803
rect 16520 21710 16593 21769
rect 16683 21710 16744 21769
rect 16520 21683 16744 21710
rect 21358 21773 21543 21792
rect 21358 21709 21412 21773
rect 21490 21709 21543 21773
rect 21358 21696 21543 21709
rect 26222 21776 26412 21792
rect 26222 21706 26264 21776
rect 26375 21706 26412 21776
rect 26222 21687 26412 21706
rect 31024 21771 31248 21792
rect 31024 21714 31080 21771
rect 31193 21714 31248 21771
rect 31024 21691 31248 21714
rect 37107 21773 37270 21793
rect 37107 21707 37146 21773
rect 37224 21707 37270 21773
rect 37107 21692 37270 21707
rect 457 21384 538 21390
rect -1736 21380 538 21384
rect -1736 21323 467 21380
rect 528 21323 538 21380
rect -1736 21317 538 21323
rect -1736 17684 -1399 21317
rect 457 21313 538 21317
rect 335 20925 559 20947
rect 335 20849 392 20925
rect 505 20849 559 20925
rect 335 20829 559 20849
rect 3808 20940 4034 20970
rect 3808 20871 3864 20940
rect 3976 20871 4034 20940
rect 3808 20844 4034 20871
rect 8623 20940 8848 20987
rect 8623 20855 8678 20940
rect 8793 20855 8848 20940
rect 8623 20822 8848 20855
rect 13856 20934 14035 20958
rect 13856 20866 13889 20934
rect 14003 20866 14035 20934
rect 13856 20835 14035 20866
rect 18231 20943 18383 20974
rect 18231 20864 18268 20943
rect 18348 20864 18383 20943
rect 18231 20834 18383 20864
rect 23408 20944 23632 20973
rect 23408 20862 23462 20944
rect 23576 20862 23632 20944
rect 23408 20832 23632 20862
rect 27831 20937 28057 20949
rect 27831 20864 27887 20937
rect 28000 20864 28057 20937
rect 27831 20833 28057 20864
rect 32984 20938 33208 20974
rect 32984 20874 33039 20938
rect 33155 20874 33208 20938
rect 32984 20848 33208 20874
rect 35736 20928 35937 20948
rect 35736 20869 35784 20928
rect 35896 20869 35937 20928
rect 35736 20845 35937 20869
rect 2128 20085 2352 20115
rect 2128 20019 2184 20085
rect 2296 20019 2352 20085
rect 2128 19995 2352 20019
rect 6832 20091 7057 20115
rect 6832 20014 6888 20091
rect 7000 20014 7057 20091
rect 6832 19995 7057 20014
rect 11704 20098 11928 20115
rect 11704 20016 11760 20098
rect 11872 20016 11928 20098
rect 11704 19995 11928 20016
rect 16540 20081 16720 20096
rect 16540 20022 16583 20081
rect 16673 20022 16720 20081
rect 16540 20004 16720 20022
rect 21355 20085 21540 20098
rect 21355 20021 21409 20085
rect 21486 20021 21540 20085
rect 21355 20006 21540 20021
rect 26228 20089 26418 20104
rect 26228 20017 26277 20089
rect 26366 20017 26418 20089
rect 26228 19999 26418 20017
rect 31023 20077 31248 20097
rect 31023 20020 31079 20077
rect 31192 20020 31248 20077
rect 31023 20003 31248 20020
rect 37092 20089 37277 20108
rect 37092 20023 37145 20089
rect 37223 20023 37277 20089
rect 37092 20006 37277 20023
rect 2128 18973 2352 19003
rect 2128 18907 2184 18973
rect 2296 18907 2352 18973
rect 2128 18883 2352 18907
rect 6832 18976 7056 19002
rect 6832 18901 6888 18976
rect 7000 18901 7056 18976
rect 6832 18883 7056 18901
rect 11704 18986 11928 19002
rect 11704 18904 11760 18986
rect 11872 18904 11928 18986
rect 11704 18883 11928 18904
rect 16540 18969 16720 18988
rect 16540 18910 16593 18969
rect 16665 18910 16720 18969
rect 16540 18896 16720 18910
rect 21371 18978 21516 18995
rect 21371 18914 21404 18978
rect 21481 18914 21516 18978
rect 21371 18897 21516 18914
rect 26221 18975 26417 18991
rect 26221 18903 26281 18975
rect 26370 18903 26417 18975
rect 26221 18887 26417 18903
rect 31024 18969 31249 18988
rect 31024 18911 31080 18969
rect 31192 18911 31249 18969
rect 31024 18894 31249 18911
rect 37099 18978 37284 18996
rect 37099 18909 37151 18978
rect 37227 18909 37284 18978
rect 37099 18894 37284 18909
rect 3807 18136 4033 18157
rect 336 18072 560 18097
rect 336 18005 392 18072
rect 505 18005 560 18072
rect 3807 18059 3863 18136
rect 3977 18059 4033 18136
rect 3807 18031 4033 18059
rect 8625 18139 8848 18176
rect 8625 18055 8680 18139
rect 8792 18055 8848 18139
rect 8625 18028 8848 18055
rect 13840 18138 14050 18175
rect 13840 18070 13888 18138
rect 14002 18070 14050 18138
rect 13840 18039 14050 18070
rect 18228 18144 18387 18174
rect 18228 18065 18269 18144
rect 18349 18065 18387 18144
rect 18228 18041 18387 18065
rect 23408 18143 23632 18167
rect 23408 18068 23464 18143
rect 23575 18068 23632 18143
rect 23408 18032 23632 18068
rect 27833 18139 28057 18167
rect 27833 18066 27889 18139
rect 28002 18066 28057 18139
rect 27833 18031 28057 18066
rect 32985 18117 33201 18139
rect 32985 18053 33038 18117
rect 33154 18053 33201 18117
rect 32985 18031 33201 18053
rect 35758 18127 35923 18147
rect 35758 18068 35784 18127
rect 35896 18068 35923 18127
rect 35758 18043 35923 18068
rect 336 17979 560 18005
rect 441 17684 524 17685
rect -1736 17675 524 17684
rect -1736 17618 451 17675
rect 514 17618 524 17675
rect -1736 17616 524 17618
rect -1736 9284 -1399 17616
rect 441 17608 524 17616
rect 2128 17300 2352 17315
rect 2128 17214 2184 17300
rect 2296 17214 2352 17300
rect 2128 17195 2352 17214
rect 6830 17291 7055 17313
rect 6830 17221 6888 17291
rect 7000 17221 7055 17291
rect 6830 17195 7055 17221
rect 11704 17282 11928 17314
rect 11704 17212 11761 17282
rect 11872 17212 11928 17282
rect 11704 17195 11928 17212
rect 16564 17278 16708 17295
rect 16564 17219 16599 17278
rect 16671 17219 16708 17278
rect 16564 17199 16708 17219
rect 21380 17285 21525 17299
rect 21380 17212 21407 17285
rect 21487 17212 21525 17285
rect 21380 17201 21525 17212
rect 26223 17285 26419 17304
rect 26223 17214 26270 17285
rect 26369 17214 26419 17285
rect 26223 17200 26419 17214
rect 31024 17279 31248 17294
rect 31024 17221 31080 17279
rect 31192 17221 31248 17279
rect 31024 17204 31248 17221
rect 37099 17289 37264 17304
rect 37099 17220 37143 17289
rect 37219 17220 37264 17289
rect 37099 17208 37264 17220
rect 2128 16181 2352 16203
rect 2128 16117 2184 16181
rect 2296 16117 2352 16181
rect 2128 16083 2352 16117
rect 6832 16173 7057 16200
rect 6832 16104 6887 16173
rect 7000 16104 7057 16173
rect 6832 16082 7057 16104
rect 11704 16180 11929 16203
rect 11704 16110 11762 16180
rect 11873 16110 11929 16180
rect 11704 16083 11929 16110
rect 16560 16175 16704 16193
rect 16560 16114 16588 16175
rect 16667 16114 16704 16175
rect 16560 16097 16704 16114
rect 21366 16181 21537 16197
rect 21366 16108 21411 16181
rect 21491 16108 21537 16181
rect 21366 16093 21537 16108
rect 26234 16176 26408 16192
rect 26234 16105 26271 16176
rect 26370 16105 26408 16176
rect 26234 16088 26408 16105
rect 31024 16171 31248 16187
rect 31024 16115 31080 16171
rect 31192 16115 31248 16171
rect 31024 16097 31248 16115
rect 37096 16175 37261 16191
rect 37096 16111 37144 16175
rect 37218 16111 37261 16175
rect 37096 16095 37261 16111
rect 335 15321 561 15359
rect 335 15254 378 15321
rect 513 15254 561 15321
rect 335 15232 561 15254
rect 3808 15332 4034 15373
rect 3808 15255 3863 15332
rect 3977 15255 4034 15332
rect 3808 15231 4034 15255
rect 8624 15343 8849 15372
rect 8624 15249 8679 15343
rect 8791 15249 8849 15343
rect 8624 15218 8849 15249
rect 13846 15338 14056 15369
rect 13846 15263 13887 15338
rect 14008 15263 14056 15338
rect 13846 15233 14056 15263
rect 18235 15336 18394 15369
rect 18235 15261 18267 15336
rect 18351 15261 18394 15336
rect 18235 15236 18394 15261
rect 23409 15324 23633 15368
rect 23409 15258 23462 15324
rect 23577 15258 23633 15324
rect 23409 15233 23633 15258
rect 27832 15334 28056 15371
rect 27832 15263 27888 15334
rect 28000 15263 28056 15334
rect 27832 15235 28056 15263
rect 32988 15339 33204 15360
rect 32988 15269 33040 15339
rect 33152 15269 33204 15339
rect 32988 15252 33204 15269
rect 35755 15333 35920 15357
rect 35755 15274 35784 15333
rect 35896 15274 35920 15333
rect 35755 15253 35920 15274
rect 2128 14495 2352 14515
rect 2128 14425 2184 14495
rect 2296 14425 2352 14495
rect 2128 14395 2352 14425
rect 6832 14489 7056 14515
rect 6832 14420 6888 14489
rect 7001 14420 7056 14489
rect 6832 14395 7056 14420
rect 11704 14494 11929 14515
rect 11704 14418 11760 14494
rect 11873 14418 11929 14494
rect 11704 14395 11929 14418
rect 16555 14478 16714 14499
rect 16555 14417 16592 14478
rect 16671 14417 16714 14478
rect 16555 14401 16714 14417
rect 21358 14481 21529 14504
rect 21358 14410 21397 14481
rect 21484 14410 21529 14481
rect 21358 14400 21529 14410
rect 26228 14483 26402 14503
rect 26228 14414 26265 14483
rect 26371 14414 26402 14483
rect 26228 14399 26402 14414
rect 31024 14479 31249 14498
rect 31024 14423 31080 14479
rect 31192 14423 31249 14479
rect 31024 14406 31249 14423
rect 37105 14489 37272 14508
rect 37105 14425 37150 14489
rect 37224 14425 37272 14489
rect 37105 14405 37272 14425
rect 2128 13383 2352 13403
rect 2128 13310 2184 13383
rect 2296 13310 2352 13383
rect 2128 13283 2352 13310
rect 6832 13374 7056 13403
rect 6832 13305 6885 13374
rect 7001 13305 7056 13374
rect 6832 13283 7056 13305
rect 11704 13384 11929 13402
rect 11704 13308 11760 13384
rect 11873 13308 11929 13384
rect 11704 13283 11929 13308
rect 16547 13372 16706 13392
rect 16547 13308 16594 13372
rect 16668 13308 16706 13372
rect 16547 13294 16706 13308
rect 21375 13376 21526 13393
rect 21375 13305 21406 13376
rect 21493 13305 21526 13376
rect 21375 13288 21526 13305
rect 26228 13380 26410 13396
rect 26228 13311 26267 13380
rect 26373 13311 26410 13380
rect 26228 13292 26410 13311
rect 31024 13370 31249 13390
rect 31024 13310 31080 13370
rect 31192 13310 31249 13370
rect 31024 13298 31249 13310
rect 37107 13376 37274 13394
rect 37107 13308 37148 13376
rect 37226 13308 37274 13376
rect 37107 13291 37274 13308
rect 3807 12535 4033 12574
rect 363 12463 532 12498
rect 363 12402 396 12463
rect 501 12402 532 12463
rect 3807 12464 3864 12535
rect 3977 12464 4033 12535
rect 3807 12432 4033 12464
rect 8624 12549 8849 12574
rect 8624 12455 8681 12549
rect 8793 12455 8849 12549
rect 8624 12429 8849 12455
rect 13830 12535 14058 12579
rect 13830 12460 13885 12535
rect 14006 12460 14058 12535
rect 13830 12432 14058 12460
rect 18216 12530 18394 12566
rect 18216 12455 18268 12530
rect 18352 12455 18394 12530
rect 18216 12431 18394 12455
rect 23408 12526 23633 12555
rect 23408 12460 23462 12526
rect 23577 12460 23633 12526
rect 23408 12432 23633 12460
rect 27833 12527 28055 12559
rect 27833 12456 27889 12527
rect 28001 12456 28055 12527
rect 27833 12431 28055 12456
rect 33004 12535 33183 12558
rect 33004 12465 33040 12535
rect 33152 12465 33183 12535
rect 33004 12445 33183 12465
rect 35750 12524 35932 12542
rect 35750 12465 35784 12524
rect 35896 12465 35932 12524
rect 35750 12442 35932 12465
rect 363 12379 532 12402
rect 2128 11700 2352 11715
rect 2128 11616 2184 11700
rect 2296 11616 2352 11700
rect 2128 11595 2352 11616
rect 6832 11684 7056 11714
rect 6832 11615 6886 11684
rect 7002 11615 7056 11684
rect 6832 11594 7056 11615
rect 11704 11686 11929 11714
rect 11704 11611 11760 11686
rect 11872 11611 11929 11686
rect 11704 11595 11929 11611
rect 16567 11681 16716 11697
rect 16567 11617 16601 11681
rect 16675 11617 16716 11681
rect 16567 11603 16716 11617
rect 21365 11686 21516 11704
rect 21365 11610 21397 11686
rect 21483 11610 21516 11686
rect 21365 11599 21516 11610
rect 26230 11687 26412 11703
rect 26230 11611 26278 11687
rect 26367 11611 26412 11687
rect 26230 11599 26412 11611
rect 31024 11685 31248 11698
rect 31024 11625 31080 11685
rect 31192 11625 31248 11685
rect 31024 11610 31248 11625
rect 37094 11686 37270 11704
rect 37094 11618 37146 11686
rect 37224 11618 37270 11686
rect 37094 11603 37270 11618
rect 2128 10581 2352 10603
rect 2128 10503 2184 10581
rect 2296 10503 2352 10581
rect 2128 10483 2352 10503
rect 6831 10576 7055 10602
rect 6831 10505 6887 10576
rect 7001 10505 7055 10576
rect 6831 10482 7055 10505
rect 11704 10583 11928 10603
rect 11704 10508 11760 10583
rect 11872 10508 11928 10583
rect 11704 10483 11928 10508
rect 16560 10574 16709 10592
rect 16560 10512 16593 10574
rect 16669 10512 16709 10574
rect 16560 10498 16709 10512
rect 21357 10576 21525 10591
rect 21357 10500 21402 10576
rect 21488 10500 21525 10576
rect 21357 10489 21525 10500
rect 26228 10582 26415 10596
rect 26228 10506 26277 10582
rect 26366 10506 26415 10582
rect 26228 10489 26415 10506
rect 31024 10574 31248 10590
rect 31024 10518 31080 10574
rect 31193 10518 31248 10574
rect 31024 10502 31248 10518
rect 37093 10579 37269 10594
rect 37093 10506 37137 10579
rect 37219 10506 37269 10579
rect 37093 10493 37269 10506
rect 336 9719 503 9744
rect 336 9654 368 9719
rect 474 9654 503 9719
rect 336 9632 503 9654
rect 3808 9741 4034 9767
rect 3808 9670 3863 9741
rect 3976 9670 4034 9741
rect 3808 9632 4034 9670
rect 8622 9730 8847 9762
rect 8622 9647 8680 9730
rect 8794 9647 8847 9730
rect 8622 9617 8847 9647
rect 13830 9735 14058 9780
rect 13830 9663 13887 9735
rect 14004 9663 14058 9735
rect 13830 9633 14058 9663
rect 18213 9735 18391 9766
rect 18213 9655 18265 9735
rect 18353 9655 18391 9735
rect 18213 9631 18391 9655
rect 23407 9726 23632 9763
rect 23407 9663 23463 9726
rect 23578 9663 23632 9726
rect 23407 9640 23632 9663
rect 27833 9733 28055 9762
rect 27833 9663 27888 9733
rect 28000 9663 28055 9733
rect 27833 9634 28055 9663
rect 33003 9732 33182 9760
rect 33003 9666 33031 9732
rect 33143 9666 33182 9732
rect 33003 9647 33182 9666
rect 35745 9732 35927 9755
rect 35745 9674 35784 9732
rect 35896 9674 35927 9732
rect 35745 9655 35927 9674
rect 334 9284 419 9288
rect -1736 9278 419 9284
rect -1736 9214 344 9278
rect 408 9214 419 9278
rect -1736 9209 419 9214
rect -1736 6631 -1399 9209
rect 334 9203 419 9209
rect 2128 8893 2352 8915
rect 2128 8813 2184 8893
rect 2296 8813 2352 8893
rect 2128 8795 2352 8813
rect 6833 8885 7057 8913
rect 6833 8814 6886 8885
rect 7000 8814 7057 8885
rect 6833 8795 7057 8814
rect 11704 8889 11928 8914
rect 11704 8811 11760 8889
rect 11872 8811 11928 8889
rect 11704 8794 11928 8811
rect 16551 8878 16727 8900
rect 16551 8816 16598 8878
rect 16674 8816 16727 8878
rect 16551 8802 16727 8816
rect 21357 8885 21525 8904
rect 21357 8811 21397 8885
rect 21484 8811 21525 8885
rect 21357 8802 21525 8811
rect 26223 8886 26410 8907
rect 26223 8811 26265 8886
rect 26364 8811 26410 8886
rect 26223 8800 26410 8811
rect 31033 8882 31231 8900
rect 31033 8826 31079 8882
rect 31192 8826 31231 8882
rect 31033 8807 31231 8826
rect 37092 8885 37270 8901
rect 37092 8812 37142 8885
rect 37224 8812 37270 8885
rect 37092 8802 37270 8812
rect 2128 7784 2352 7803
rect 2128 7714 2184 7784
rect 2296 7714 2352 7784
rect 2128 7683 2352 7714
rect 6832 7773 7056 7802
rect 6832 7708 6888 7773
rect 7000 7708 7056 7773
rect 6832 7684 7056 7708
rect 11704 7781 11928 7802
rect 11704 7703 11760 7781
rect 11872 7703 11928 7781
rect 11704 7683 11928 7703
rect 16540 7772 16716 7791
rect 16540 7706 16589 7772
rect 16670 7706 16716 7772
rect 16540 7693 16716 7706
rect 21363 7779 21532 7793
rect 21363 7705 21404 7779
rect 21491 7705 21532 7779
rect 21363 7689 21532 7705
rect 26231 7783 26414 7796
rect 26231 7708 26273 7783
rect 26372 7708 26414 7783
rect 26231 7693 26414 7708
rect 31031 7772 31229 7790
rect 31031 7716 31079 7772
rect 31192 7716 31229 7772
rect 31031 7697 31229 7716
rect 37097 7779 37275 7794
rect 37097 7711 37144 7779
rect 37228 7711 37275 7779
rect 37097 7695 37275 7711
rect 3807 6935 4033 6967
rect 337 6874 561 6900
rect 337 6805 390 6874
rect 505 6805 561 6874
rect 3807 6854 3863 6935
rect 3977 6854 4033 6935
rect 3807 6832 4033 6854
rect 8623 6928 8848 6965
rect 8623 6849 8679 6928
rect 8791 6849 8848 6928
rect 8623 6824 8848 6849
rect 13832 6938 14058 6973
rect 13832 6866 13886 6938
rect 14003 6866 14058 6938
rect 13832 6838 14058 6866
rect 18225 6956 18392 6977
rect 18225 6876 18263 6956
rect 18351 6876 18392 6956
rect 18225 6855 18392 6876
rect 23406 6928 23634 6962
rect 23406 6865 23462 6928
rect 23577 6865 23634 6928
rect 23406 6834 23634 6865
rect 27831 6939 28053 6967
rect 27831 6869 27887 6939
rect 27999 6869 28053 6939
rect 27831 6832 28053 6869
rect 33009 6930 33190 6951
rect 33009 6864 33041 6930
rect 33153 6864 33190 6930
rect 33009 6842 33190 6864
rect 35737 6921 35937 6945
rect 35737 6863 35784 6921
rect 35896 6863 35937 6921
rect 35737 6839 35937 6863
rect 337 6779 561 6805
rect -1736 6559 621 6631
rect -1736 3684 -1399 6559
rect 549 6489 621 6559
rect 544 6479 628 6489
rect 544 6416 554 6479
rect 618 6416 628 6479
rect 544 6406 628 6416
rect 2128 6088 2352 6115
rect 2128 6012 2184 6088
rect 2296 6012 2352 6088
rect 2128 5995 2352 6012
rect 6832 6081 7056 6115
rect 6832 6016 6888 6081
rect 7000 6016 7056 6081
rect 6832 5995 7056 6016
rect 11703 6089 11927 6114
rect 11703 6016 11761 6089
rect 11874 6016 11927 6089
rect 11703 5995 11927 6016
rect 16558 6082 16730 6104
rect 16558 6016 16593 6082
rect 16674 6016 16730 6082
rect 16558 5998 16730 6016
rect 21359 6083 21528 6105
rect 21359 6011 21400 6083
rect 21485 6011 21528 6083
rect 21359 6001 21528 6011
rect 26232 6090 26415 6102
rect 26232 6010 26275 6090
rect 26367 6010 26415 6090
rect 26232 5999 26415 6010
rect 31049 6082 31220 6098
rect 31049 6026 31080 6082
rect 31193 6026 31220 6082
rect 31049 6009 31220 6026
rect 37090 6083 37270 6101
rect 37090 6015 37140 6083
rect 37224 6015 37270 6083
rect 37090 6002 37270 6015
rect 2128 4984 2353 5003
rect 2128 4910 2184 4984
rect 2296 4910 2353 4984
rect 2128 4883 2353 4910
rect 6832 4974 7056 5003
rect 6832 4903 6888 4974
rect 7001 4903 7056 4974
rect 6832 4883 7056 4903
rect 11704 4980 11929 5002
rect 11704 4907 11759 4980
rect 11872 4907 11929 4980
rect 11704 4883 11929 4907
rect 16545 4976 16717 4993
rect 16545 4906 16589 4976
rect 16672 4906 16717 4976
rect 16545 4887 16717 4906
rect 21375 4974 21532 4993
rect 21375 4902 21408 4974
rect 21493 4902 21532 4974
rect 21375 4887 21532 4902
rect 26242 4980 26415 4996
rect 26242 4900 26281 4980
rect 26373 4900 26415 4980
rect 31050 4977 31221 4990
rect 31050 4921 31080 4977
rect 31192 4921 31221 4977
rect 31050 4901 31221 4921
rect 37100 4976 37280 4992
rect 37100 4910 37140 4976
rect 37228 4910 37280 4976
rect 26242 4886 26415 4900
rect 37100 4893 37280 4910
rect 336 4141 561 4200
rect 336 4062 390 4141
rect 507 4062 561 4141
rect 336 4028 561 4062
rect 3808 4139 4032 4172
rect 3808 4058 3863 4139
rect 3977 4058 4032 4139
rect 3808 4031 4032 4058
rect 8624 4129 8849 4164
rect 8624 4052 8680 4129
rect 8793 4052 8849 4129
rect 8624 4025 8849 4052
rect 13831 4135 14057 4166
rect 13831 4060 13887 4135
rect 14000 4060 14057 4135
rect 13831 4033 14057 4060
rect 18222 4141 18389 4170
rect 18222 4066 18267 4141
rect 18360 4066 18389 4141
rect 18222 4048 18389 4066
rect 23407 4127 23635 4161
rect 23407 4056 23460 4127
rect 23576 4056 23635 4127
rect 23407 4033 23635 4056
rect 27834 4123 28056 4160
rect 27834 4050 27887 4123
rect 28001 4050 28056 4123
rect 27834 4025 28056 4050
rect 32997 4136 33178 4158
rect 32997 4072 33030 4136
rect 33139 4072 33178 4136
rect 32997 4049 33178 4072
rect 35742 4130 35942 4159
rect 35742 4074 35783 4130
rect 35896 4074 35942 4130
rect 35742 4053 35942 4074
rect 318 3684 401 3687
rect -1736 3677 401 3684
rect -1736 3617 328 3677
rect 391 3617 401 3677
rect -1736 3614 401 3617
rect -1736 2800 -1399 3614
rect 318 3607 401 3614
rect 2128 3293 2352 3315
rect 2128 3214 2184 3293
rect 2296 3214 2352 3293
rect 2128 3195 2352 3214
rect 6832 3288 7056 3314
rect 6832 3217 6888 3288
rect 7001 3217 7056 3288
rect 6832 3194 7056 3217
rect 11701 3284 11926 3314
rect 11701 3209 11757 3284
rect 11875 3209 11926 3284
rect 11701 3195 11926 3209
rect 16560 3288 16719 3302
rect 16560 3218 16594 3288
rect 16677 3218 16719 3288
rect 16560 3202 16719 3218
rect 21371 3283 21528 3303
rect 21371 3212 21401 3283
rect 21486 3212 21528 3283
rect 21371 3197 21528 3212
rect 26229 3290 26402 3309
rect 26229 3210 26264 3290
rect 26360 3210 26402 3290
rect 26229 3199 26402 3210
rect 31051 3278 31233 3299
rect 31051 3222 31080 3278
rect 31192 3222 31233 3278
rect 31051 3204 31233 3222
rect 37093 3285 37278 3305
rect 37093 3219 37137 3285
rect 37225 3219 37278 3285
rect 37093 3206 37278 3219
rect 2128 2172 2352 2203
rect 2128 2104 2184 2172
rect 2296 2104 2352 2172
rect 2128 2083 2352 2104
rect 6832 2173 7056 2204
rect 6832 2104 6887 2173
rect 7001 2104 7056 2173
rect 6832 2084 7056 2104
rect 11702 2181 11929 2200
rect 11702 2106 11758 2181
rect 11876 2106 11929 2181
rect 11702 2085 11929 2106
rect 16553 2177 16712 2194
rect 16553 2104 16595 2177
rect 16675 2104 16712 2177
rect 16553 2094 16712 2104
rect 21376 2174 21524 2196
rect 21376 2103 21403 2174
rect 21488 2103 21524 2174
rect 21376 2084 21524 2103
rect 26227 2179 26412 2195
rect 26227 2099 26276 2179
rect 26372 2099 26412 2179
rect 31046 2178 31228 2194
rect 31046 2117 31079 2178
rect 31193 2117 31228 2178
rect 31046 2099 31228 2117
rect 26227 2088 26412 2099
rect 3808 1332 4032 1378
rect 3808 1265 3864 1332
rect 3976 1265 4032 1332
rect 3808 1232 4032 1265
rect 8625 1334 8849 1364
rect 8625 1257 8679 1334
rect 8792 1257 8849 1334
rect 8625 1231 8849 1257
rect 13834 1328 14055 1363
rect 13834 1255 13872 1328
rect 14002 1255 14055 1328
rect 13834 1219 14055 1255
rect 18198 1335 18424 1361
rect 18198 1260 18262 1335
rect 18355 1260 18424 1335
rect 18198 1233 18424 1260
rect 23409 1342 23632 1368
rect 23409 1271 23462 1342
rect 23578 1271 23632 1342
rect 23409 1233 23632 1271
rect 27832 1330 28059 1357
rect 27832 1257 27887 1330
rect 28001 1257 28059 1330
rect 27832 1233 28059 1257
rect 33008 1329 33186 1356
rect 33008 1265 33043 1329
rect 33152 1265 33186 1329
rect 33008 1241 33186 1265
rect 2128 489 2352 515
rect 2128 416 2184 489
rect 2296 416 2352 489
rect 2128 395 2352 416
rect 6831 487 7057 515
rect 6831 418 6887 487
rect 7001 418 7057 487
rect 6831 395 7057 418
rect 11704 487 11931 511
rect 11704 410 11760 487
rect 11872 410 11931 487
rect 11704 396 11931 410
rect 16529 485 16723 502
rect 16529 412 16588 485
rect 16668 412 16723 485
rect 16529 401 16723 412
rect 21369 480 21517 507
rect 21369 408 21402 480
rect 21481 408 21517 480
rect 21369 395 21517 408
rect 26229 483 26414 505
rect 26229 406 26275 483
rect 26363 406 26414 483
rect 26229 398 26414 406
rect 31041 482 31228 504
rect 31041 421 31079 482
rect 31193 421 31228 482
rect 31041 402 31228 421
<< via3 >>
rect 35783 26137 35896 26199
rect 37139 25335 37230 25411
rect 35784 25176 35897 25238
rect 37137 24378 37228 24454
rect 391 22657 504 22733
rect 8680 23169 8793 23243
rect 13888 23184 13944 23240
rect 18283 23184 18339 23240
rect 23493 23184 23549 23240
rect 27862 23179 28000 23251
rect 35784 24221 35896 24283
rect 37140 23426 37220 23495
rect 35784 23238 35896 23300
rect 3881 22614 3971 22672
rect 11761 22389 11874 22465
rect 16605 22400 16661 22456
rect 21421 22400 21477 22456
rect 26292 22400 26348 22456
rect 31111 22400 31167 22456
rect 37137 22449 37216 22518
rect 37216 22449 37217 22518
rect 2184 21703 2296 21777
rect 6887 21698 7001 21776
rect 11760 21700 11873 21782
rect 16593 21710 16683 21769
rect 21412 21709 21490 21773
rect 26264 21706 26375 21776
rect 31080 21714 31193 21771
rect 37146 21707 37224 21773
rect 392 20849 505 20925
rect 3864 20871 3976 20940
rect 8678 20855 8793 20940
rect 13889 20866 14003 20934
rect 18268 20864 18348 20943
rect 23462 20862 23576 20944
rect 27887 20864 28000 20937
rect 33039 20874 33155 20938
rect 35784 20869 35896 20928
rect 2184 20019 2296 20085
rect 6888 20014 7000 20091
rect 11760 20016 11872 20098
rect 16583 20022 16673 20081
rect 21409 20021 21486 20085
rect 26277 20017 26366 20089
rect 31079 20020 31192 20077
rect 37145 20023 37223 20089
rect 2184 18907 2296 18973
rect 6888 18901 7000 18976
rect 11760 18904 11872 18986
rect 16593 18910 16665 18969
rect 21404 18914 21481 18978
rect 26281 18903 26370 18975
rect 31080 18911 31192 18969
rect 37151 18909 37227 18978
rect 392 18005 505 18072
rect 3863 18059 3977 18136
rect 8680 18055 8792 18139
rect 13888 18070 14002 18138
rect 18269 18065 18349 18144
rect 23464 18068 23575 18143
rect 27889 18066 28002 18139
rect 33038 18053 33154 18117
rect 35784 18068 35896 18127
rect 2184 17214 2296 17300
rect 6888 17221 7000 17291
rect 11761 17212 11872 17282
rect 16599 17219 16671 17278
rect 21407 17212 21487 17285
rect 26270 17214 26369 17285
rect 31080 17221 31192 17279
rect 37143 17220 37219 17289
rect 2184 16117 2296 16181
rect 6887 16104 7000 16173
rect 11762 16110 11873 16180
rect 16588 16114 16667 16175
rect 21411 16108 21491 16181
rect 26271 16105 26370 16176
rect 31080 16115 31192 16171
rect 37144 16111 37218 16175
rect 378 15254 513 15321
rect 3863 15255 3977 15332
rect 8679 15249 8791 15343
rect 13887 15263 14008 15338
rect 18267 15261 18351 15336
rect 23462 15258 23577 15324
rect 33040 15269 33152 15339
rect 35784 15274 35896 15333
rect 2184 14425 2296 14495
rect 6888 14420 7001 14489
rect 11760 14418 11873 14494
rect 16592 14417 16671 14478
rect 21397 14410 21484 14481
rect 26265 14414 26371 14483
rect 31080 14423 31192 14479
rect 37150 14425 37224 14489
rect 2184 13310 2296 13383
rect 6885 13305 7001 13374
rect 11760 13308 11873 13384
rect 16594 13308 16668 13372
rect 21406 13305 21493 13376
rect 26267 13311 26373 13380
rect 31080 13310 31192 13370
rect 37148 13308 37226 13376
rect 396 12402 501 12463
rect 3864 12464 3977 12535
rect 8681 12455 8793 12549
rect 13885 12460 14006 12535
rect 18268 12455 18352 12530
rect 23462 12460 23577 12526
rect 27889 12456 28001 12527
rect 33040 12465 33152 12535
rect 35784 12465 35896 12524
rect 2184 11616 2296 11700
rect 6886 11615 7002 11684
rect 11760 11611 11872 11686
rect 16601 11617 16675 11681
rect 21397 11610 21483 11686
rect 26278 11611 26367 11687
rect 31080 11625 31192 11685
rect 37146 11618 37224 11686
rect 2184 10503 2296 10581
rect 6887 10505 7001 10576
rect 11760 10508 11872 10583
rect 16593 10512 16669 10574
rect 21402 10500 21488 10576
rect 26277 10506 26366 10582
rect 31080 10518 31193 10574
rect 37137 10506 37219 10579
rect 368 9654 474 9719
rect 3863 9670 3976 9741
rect 8680 9647 8794 9730
rect 13887 9663 14004 9735
rect 18265 9655 18353 9735
rect 23463 9663 23578 9726
rect 27888 9663 28000 9733
rect 33031 9666 33143 9732
rect 35784 9674 35896 9732
rect 2184 8813 2296 8893
rect 6886 8814 7000 8885
rect 11760 8811 11872 8889
rect 16598 8816 16674 8878
rect 21397 8811 21484 8885
rect 26265 8811 26364 8886
rect 31079 8826 31192 8882
rect 37142 8812 37224 8885
rect 2184 7714 2296 7784
rect 6888 7708 7000 7773
rect 11760 7703 11872 7781
rect 16589 7706 16670 7772
rect 21404 7705 21491 7779
rect 26273 7708 26372 7783
rect 31079 7716 31192 7772
rect 37144 7711 37228 7779
rect 390 6805 505 6874
rect 3863 6854 3977 6935
rect 8679 6849 8791 6928
rect 13886 6866 14003 6938
rect 18263 6876 18351 6956
rect 23462 6865 23577 6928
rect 33041 6864 33153 6930
rect 35784 6863 35896 6921
rect 2184 6012 2296 6088
rect 6888 6016 7000 6081
rect 11761 6016 11874 6089
rect 16593 6016 16674 6082
rect 21400 6011 21485 6083
rect 26275 6010 26367 6090
rect 31080 6026 31193 6082
rect 37140 6015 37224 6083
rect 2184 4910 2296 4984
rect 6888 4903 7001 4974
rect 11759 4907 11872 4980
rect 16589 4906 16672 4976
rect 21408 4902 21493 4974
rect 26281 4900 26373 4980
rect 31080 4921 31192 4977
rect 37140 4910 37228 4976
rect 390 4062 507 4141
rect 3863 4058 3977 4139
rect 8680 4052 8793 4129
rect 13887 4060 14000 4135
rect 18267 4066 18360 4141
rect 23460 4056 23576 4127
rect 27887 4050 28001 4123
rect 33030 4072 33139 4136
rect 35783 4074 35896 4130
rect 2184 3214 2296 3293
rect 6888 3217 7001 3288
rect 11757 3209 11875 3284
rect 16594 3218 16677 3288
rect 21401 3212 21486 3283
rect 26264 3210 26360 3290
rect 31080 3222 31192 3278
rect 37137 3219 37225 3285
rect 2184 2104 2296 2172
rect 6887 2104 7001 2173
rect 11758 2106 11876 2181
rect 16595 2104 16675 2177
rect 21403 2103 21488 2174
rect 26276 2099 26372 2179
rect 31079 2117 31193 2178
rect 3864 1265 3976 1332
rect 8679 1257 8792 1334
rect 13872 1255 14002 1328
rect 18262 1260 18355 1335
rect 23462 1271 23578 1342
rect 27887 1257 28001 1330
rect 33043 1265 33152 1329
rect 2184 416 2296 489
rect 6887 418 7001 487
rect 11760 410 11872 487
rect 16588 412 16668 485
rect 21402 408 21481 480
rect 26275 406 26363 483
rect 31079 421 31193 482
<< metal4 >>
rect -6209 30193 -854 30196
rect -6209 30190 44816 30193
rect -6209 29717 46985 30190
rect -6209 27719 46986 29717
rect -6209 27715 -854 27719
rect -6204 20317 -3615 27715
rect 280 22733 616 27719
rect 280 22657 391 22733
rect 504 22657 616 22733
rect 280 22260 616 22657
rect 311 22120 616 22260
rect 280 21516 616 22120
rect 3752 22672 4088 27719
rect 3752 22614 3881 22672
rect 3971 22614 4088 22672
rect 336 21366 616 21516
rect -6204 20293 -5232 20317
rect -4434 20293 -3615 20317
rect -6204 19920 -5297 20293
rect -4423 19920 -3615 20293
rect -6204 19913 -5232 19920
rect -4434 19913 -3615 19920
rect -6204 17438 -3615 19913
rect -6204 17031 -5228 17438
rect -4377 17031 -3615 17438
rect -6204 14586 -3615 17031
rect -6204 14179 -5317 14586
rect -4466 14179 -3615 14586
rect -6204 11850 -3615 14179
rect -6204 11443 -5253 11850
rect -4402 11443 -3615 11850
rect -6204 9046 -3615 11443
rect -6204 8639 -5326 9046
rect -4475 8639 -3615 9046
rect -6204 6309 -3615 8639
rect -6204 5902 -5235 6309
rect -4384 5902 -3615 6309
rect -6204 3505 -3615 5902
rect -6204 3098 -5349 3505
rect -4498 3098 -3615 3505
rect -6204 653 -3615 3098
rect 280 20925 616 21366
rect 280 20849 392 20925
rect 505 20849 616 20925
rect 280 20145 616 20849
rect 280 20027 364 20145
rect 530 20027 616 20145
rect 280 18072 616 20027
rect 280 18005 392 18072
rect 505 18005 616 18072
rect 280 17298 616 18005
rect 280 17180 359 17298
rect 525 17180 616 17298
rect 280 15321 616 17180
rect 280 15254 378 15321
rect 513 15254 616 15321
rect 280 14428 616 15254
rect 280 14310 362 14428
rect 528 14310 616 14428
rect 280 12463 616 14310
rect 280 12402 396 12463
rect 501 12402 616 12463
rect 280 11709 616 12402
rect 280 11591 365 11709
rect 531 11591 616 11709
rect 280 9719 616 11591
rect 280 9654 368 9719
rect 474 9654 616 9719
rect 280 8901 616 9654
rect 280 8783 369 8901
rect 535 8783 616 8901
rect 280 6874 616 8783
rect 280 6805 390 6874
rect 505 6805 616 6874
rect 280 6151 616 6805
rect 280 6033 370 6151
rect 536 6033 616 6151
rect 280 4141 616 6033
rect 280 4062 390 4141
rect 507 4062 616 4141
rect 280 3352 616 4062
rect 280 3234 364 3352
rect 530 3234 616 3352
rect 280 699 616 3234
rect 2072 21788 2408 22014
rect 2072 21693 2169 21788
rect 2306 21693 2408 21788
rect 2072 20085 2408 21693
rect 2072 20019 2184 20085
rect 2296 20019 2408 20085
rect 2072 18988 2408 20019
rect 2072 18893 2169 18988
rect 2306 18893 2408 18988
rect 2072 17300 2408 18893
rect 2072 17214 2184 17300
rect 2296 17214 2408 17300
rect 2072 16197 2408 17214
rect 2072 16102 2171 16197
rect 2308 16102 2408 16197
rect 2072 14495 2408 16102
rect 2072 14425 2184 14495
rect 2296 14425 2408 14495
rect 2072 13393 2408 14425
rect 2072 13298 2175 13393
rect 2312 13298 2408 13393
rect 2072 11700 2408 13298
rect 2072 11616 2184 11700
rect 2296 11616 2408 11700
rect 2072 10591 2408 11616
rect 2072 10496 2172 10591
rect 2309 10496 2408 10591
rect 2072 8893 2408 10496
rect 2072 8813 2184 8893
rect 2296 8813 2408 8893
rect 2072 7795 2408 8813
rect 2072 7700 2170 7795
rect 2307 7700 2408 7795
rect 2072 6088 2408 7700
rect 2072 6012 2184 6088
rect 2296 6012 2408 6088
rect 2072 4995 2408 6012
rect 2072 4900 2173 4995
rect 2310 4900 2408 4995
rect 2072 3293 2408 4900
rect 2072 3214 2184 3293
rect 2296 3214 2408 3293
rect 2072 2187 2408 3214
rect 2072 2092 2171 2187
rect 2308 2092 2408 2187
rect -6204 246 -5047 653
rect -4196 246 -3615 653
rect -6204 -1009 -3615 246
rect 275 489 617 699
rect 275 371 359 489
rect 525 371 617 489
rect 275 -1002 617 371
rect 2072 489 2408 2092
rect 2072 416 2184 489
rect 2296 416 2408 489
rect 2072 305 2408 416
rect 2069 168 2408 305
rect 3752 20940 4088 22614
rect 8568 23243 8904 27719
rect 8568 23169 8680 23243
rect 8793 23169 8904 23243
rect 3752 20871 3864 20940
rect 3976 20871 4088 20940
rect 3752 20139 4088 20871
rect 3752 20021 3835 20139
rect 4001 20021 4088 20139
rect 3752 18136 4088 20021
rect 3752 18059 3863 18136
rect 3977 18059 4088 18136
rect 3752 17282 4088 18059
rect 3752 17164 3826 17282
rect 3992 17164 4088 17282
rect 3752 15332 4088 17164
rect 3752 15255 3863 15332
rect 3977 15255 4088 15332
rect 3752 14441 4088 15255
rect 3752 14323 3830 14441
rect 3996 14323 4088 14441
rect 3752 12535 4088 14323
rect 3752 12464 3864 12535
rect 3977 12464 4088 12535
rect 3752 11708 4088 12464
rect 3752 11590 3841 11708
rect 4007 11590 4088 11708
rect 3752 9741 4088 11590
rect 3752 9670 3863 9741
rect 3976 9670 4088 9741
rect 3752 8887 4088 9670
rect 3752 8769 3834 8887
rect 4000 8769 4088 8887
rect 3752 6935 4088 8769
rect 3752 6854 3863 6935
rect 3977 6854 4088 6935
rect 3752 6141 4088 6854
rect 3752 6023 3825 6141
rect 3991 6023 4088 6141
rect 3752 4139 4088 6023
rect 3752 4058 3863 4139
rect 3977 4058 4088 4139
rect 3752 3339 4088 4058
rect 3752 3221 3837 3339
rect 4003 3221 4088 3339
rect 3752 1332 4088 3221
rect 3752 1265 3864 1332
rect 3976 1265 4088 1332
rect 3752 502 4088 1265
rect 3752 384 3831 502
rect 3997 384 4088 502
rect 3752 230 4088 384
rect 3751 168 4088 230
rect 6776 21787 7112 22004
rect 6776 21692 6877 21787
rect 7014 21692 7112 21787
rect 6776 20091 7112 21692
rect 6776 20014 6888 20091
rect 7000 20014 7112 20091
rect 6776 18988 7112 20014
rect 6776 18893 6875 18988
rect 7012 18893 7112 18988
rect 6776 17291 7112 18893
rect 6776 17221 6888 17291
rect 7000 17221 7112 17291
rect 6776 16186 7112 17221
rect 6776 16091 6873 16186
rect 7010 16091 7112 16186
rect 6776 14489 7112 16091
rect 6776 14420 6888 14489
rect 7001 14420 7112 14489
rect 6776 13388 7112 14420
rect 6776 13293 6871 13388
rect 7008 13293 7112 13388
rect 6776 11684 7112 13293
rect 6776 11615 6886 11684
rect 7002 11615 7112 11684
rect 6776 10592 7112 11615
rect 6776 10497 6876 10592
rect 7013 10497 7112 10592
rect 6776 8885 7112 10497
rect 6776 8814 6886 8885
rect 7000 8814 7112 8885
rect 6776 7787 7112 8814
rect 6776 7692 6872 7787
rect 7009 7692 7112 7787
rect 6776 6081 7112 7692
rect 6776 6016 6888 6081
rect 7000 6016 7112 6081
rect 6776 4990 7112 6016
rect 6776 4895 6872 4990
rect 7009 4895 7112 4990
rect 6776 3288 7112 4895
rect 6776 3217 6888 3288
rect 7001 3217 7112 3288
rect 6776 2190 7112 3217
rect 6776 2095 6874 2190
rect 7011 2095 7112 2190
rect 6776 487 7112 2095
rect 6776 418 6887 487
rect 7001 418 7112 487
rect 2069 -252 2406 168
rect 2069 -402 2404 -252
rect 2069 -657 2128 -402
rect 2367 -657 2404 -402
rect 2069 -711 2404 -657
rect 3751 -1002 4085 168
rect 6776 0 7112 418
rect 8568 20940 8904 23169
rect 13776 23240 14112 27719
rect 13776 23184 13888 23240
rect 13944 23184 14112 23240
rect 8568 20855 8678 20940
rect 8793 20855 8904 20940
rect 8568 20161 8904 20855
rect 8568 20043 8650 20161
rect 8816 20043 8904 20161
rect 8568 18139 8904 20043
rect 8568 18055 8680 18139
rect 8792 18055 8904 18139
rect 8568 17284 8904 18055
rect 8568 17166 8652 17284
rect 8818 17166 8904 17284
rect 8568 15343 8904 17166
rect 8568 15249 8679 15343
rect 8791 15249 8904 15343
rect 8568 14437 8904 15249
rect 8568 14319 8642 14437
rect 8808 14319 8904 14437
rect 8568 12549 8904 14319
rect 8568 12455 8681 12549
rect 8793 12455 8904 12549
rect 8568 11696 8904 12455
rect 8568 11578 8663 11696
rect 8829 11578 8904 11696
rect 8568 9730 8904 11578
rect 8568 9647 8680 9730
rect 8794 9647 8904 9730
rect 8568 8887 8904 9647
rect 8568 8769 8649 8887
rect 8815 8769 8904 8887
rect 8568 6928 8904 8769
rect 8568 6849 8679 6928
rect 8791 6849 8904 6928
rect 8568 6137 8904 6849
rect 8568 6019 8664 6137
rect 8830 6019 8904 6137
rect 8568 4129 8904 6019
rect 8568 4052 8680 4129
rect 8793 4052 8904 4129
rect 8568 3357 8904 4052
rect 8568 3239 8657 3357
rect 8823 3239 8904 3357
rect 8568 1334 8904 3239
rect 8568 1257 8679 1334
rect 8792 1257 8904 1334
rect 8568 483 8904 1257
rect 8568 365 8648 483
rect 8814 365 8904 483
rect 8568 56 8904 365
rect 11648 22465 11984 22996
rect 11648 22389 11761 22465
rect 11874 22389 11984 22465
rect 11648 21791 11984 22389
rect 11648 21696 11750 21791
rect 11887 21696 11984 21791
rect 11648 20098 11984 21696
rect 11648 20016 11760 20098
rect 11872 20016 11984 20098
rect 11648 18989 11984 20016
rect 11648 18894 11745 18989
rect 11882 18894 11984 18989
rect 11648 17282 11984 18894
rect 11648 17212 11761 17282
rect 11872 17212 11984 17282
rect 11648 16192 11984 17212
rect 11648 16097 11748 16192
rect 11885 16097 11984 16192
rect 11648 14494 11984 16097
rect 11648 14418 11760 14494
rect 11873 14418 11984 14494
rect 11648 13394 11984 14418
rect 11648 13299 11743 13394
rect 11880 13299 11984 13394
rect 11648 11686 11984 13299
rect 11648 11611 11760 11686
rect 11872 11611 11984 11686
rect 11648 10589 11984 11611
rect 11648 10494 11745 10589
rect 11882 10494 11984 10589
rect 11648 8889 11984 10494
rect 11648 8811 11760 8889
rect 11872 8811 11984 8889
rect 11648 7789 11984 8811
rect 11648 7694 11746 7789
rect 11883 7694 11984 7789
rect 11648 6089 11984 7694
rect 11648 6016 11761 6089
rect 11874 6016 11984 6089
rect 11648 4991 11984 6016
rect 11648 4896 11745 4991
rect 11882 4896 11984 4991
rect 11648 3284 11984 4896
rect 11648 3209 11757 3284
rect 11875 3209 11984 3284
rect 11648 2191 11984 3209
rect 13776 20934 14112 23184
rect 18144 24528 18480 27719
rect 18144 23240 18481 24528
rect 18144 23184 18283 23240
rect 18339 23184 18481 23240
rect 13776 20866 13889 20934
rect 14003 20866 14112 20934
rect 13776 20137 14112 20866
rect 13776 20019 13853 20137
rect 14019 20019 14112 20137
rect 13776 18138 14112 20019
rect 13776 18070 13888 18138
rect 14002 18070 14112 18138
rect 13776 17293 14112 18070
rect 13776 17175 13849 17293
rect 14015 17175 14112 17293
rect 13776 15338 14112 17175
rect 13776 15263 13887 15338
rect 14008 15263 14112 15338
rect 13776 14426 14112 15263
rect 13776 14308 13851 14426
rect 14017 14308 14112 14426
rect 13776 12535 14112 14308
rect 13776 12460 13885 12535
rect 14006 12460 14112 12535
rect 13776 11723 14112 12460
rect 13776 11605 13858 11723
rect 14024 11605 14112 11723
rect 13776 9735 14112 11605
rect 13776 9663 13887 9735
rect 14004 9663 14112 9735
rect 13776 8891 14112 9663
rect 13776 8773 13869 8891
rect 14035 8773 14112 8891
rect 13776 6938 14112 8773
rect 13776 6866 13886 6938
rect 14003 6866 14112 6938
rect 13776 6132 14112 6866
rect 13776 6014 13856 6132
rect 14022 6014 14112 6132
rect 13776 4135 14112 6014
rect 13776 4060 13887 4135
rect 14000 4060 14112 4135
rect 13776 3354 14112 4060
rect 13776 3236 13858 3354
rect 14024 3236 14112 3354
rect 13776 2440 14112 3236
rect 16464 22456 16800 22700
rect 16464 22400 16605 22456
rect 16661 22400 16800 22456
rect 16464 21791 16800 22400
rect 16464 21696 16568 21791
rect 16705 21696 16800 21791
rect 16464 20081 16800 21696
rect 16464 20022 16583 20081
rect 16673 20022 16800 20081
rect 16464 18989 16800 20022
rect 16464 18894 16563 18989
rect 16700 18894 16800 18989
rect 16464 17278 16800 18894
rect 16464 17219 16599 17278
rect 16671 17219 16800 17278
rect 16464 16194 16800 17219
rect 16464 16099 16561 16194
rect 16698 16099 16800 16194
rect 16464 14478 16800 16099
rect 16464 14417 16592 14478
rect 16671 14417 16800 14478
rect 16464 13393 16800 14417
rect 16464 13298 16562 13393
rect 16699 13298 16800 13393
rect 16464 11681 16800 13298
rect 16464 11617 16601 11681
rect 16675 11617 16800 11681
rect 16464 10594 16800 11617
rect 16464 10499 16565 10594
rect 16702 10499 16800 10594
rect 16464 8878 16800 10499
rect 16464 8816 16598 8878
rect 16674 8816 16800 8878
rect 16464 7790 16800 8816
rect 16464 7695 16561 7790
rect 16698 7695 16800 7790
rect 16464 6082 16800 7695
rect 16464 6016 16593 6082
rect 16674 6016 16800 6082
rect 16464 4984 16800 6016
rect 16464 4889 16561 4984
rect 16698 4889 16800 4984
rect 16464 3288 16800 4889
rect 16464 3218 16594 3288
rect 16677 3218 16800 3288
rect 11648 2096 11748 2191
rect 11885 2096 11984 2191
rect 11648 487 11984 2096
rect 11648 410 11760 487
rect 11872 410 11984 487
rect 11648 174 11984 410
rect 6778 -101 7112 0
rect 6778 -252 7113 -101
rect 6779 -431 7113 -252
rect 6779 -696 6823 -431
rect 7082 -696 7113 -431
rect 6779 -745 7113 -696
rect 8570 -1002 8904 56
rect 11643 0 11984 174
rect 13775 1328 14114 2440
rect 13775 1255 13872 1328
rect 14002 1255 14114 1328
rect 13775 484 14114 1255
rect 13775 366 13863 484
rect 14029 366 14114 484
rect 11643 -252 11982 0
rect 11643 -393 11981 -252
rect 11643 -606 11709 -393
rect 11938 -606 11981 -393
rect 11643 -748 11981 -606
rect 13775 -1002 14114 366
rect 16464 2190 16800 3218
rect 16464 2095 16565 2190
rect 16702 2095 16800 2190
rect 16464 485 16800 2095
rect 16464 412 16588 485
rect 16668 412 16800 485
rect 16464 56 16800 412
rect 16466 -252 16800 56
rect 18144 20943 18481 23184
rect 23352 23240 23688 27719
rect 23352 23184 23493 23240
rect 23549 23184 23688 23240
rect 18144 20864 18268 20943
rect 18348 20864 18481 20943
rect 18144 20142 18481 20864
rect 18144 20024 18229 20142
rect 18395 20024 18481 20142
rect 18144 18144 18481 20024
rect 18144 18065 18269 18144
rect 18349 18065 18481 18144
rect 18144 17275 18481 18065
rect 18144 17157 18202 17275
rect 18368 17157 18481 17275
rect 18144 15336 18481 17157
rect 18144 15261 18267 15336
rect 18351 15261 18481 15336
rect 18144 14433 18481 15261
rect 18144 14315 18237 14433
rect 18403 14315 18481 14433
rect 18144 12530 18481 14315
rect 18144 12455 18268 12530
rect 18352 12455 18481 12530
rect 18144 11689 18481 12455
rect 18144 11571 18236 11689
rect 18402 11571 18481 11689
rect 18144 9735 18481 11571
rect 18144 9655 18265 9735
rect 18353 9655 18481 9735
rect 18144 8891 18481 9655
rect 18144 8773 18240 8891
rect 18406 8773 18481 8891
rect 18144 6956 18481 8773
rect 18144 6876 18263 6956
rect 18351 6876 18481 6956
rect 18144 6146 18481 6876
rect 18144 6028 18232 6146
rect 18398 6028 18481 6146
rect 18144 4141 18481 6028
rect 18144 4066 18267 4141
rect 18360 4066 18481 4141
rect 18144 3358 18481 4066
rect 18144 3240 18226 3358
rect 18392 3240 18481 3358
rect 18144 1335 18481 3240
rect 18144 1260 18262 1335
rect 18355 1260 18481 1335
rect 18144 499 18481 1260
rect 18144 381 18221 499
rect 18387 381 18481 499
rect 18144 123 18481 381
rect 21280 22456 21616 22791
rect 21280 22400 21421 22456
rect 21477 22400 21616 22456
rect 21280 21788 21616 22400
rect 21280 21693 21386 21788
rect 21523 21693 21616 21788
rect 21280 20085 21616 21693
rect 21280 20021 21409 20085
rect 21486 20021 21616 20085
rect 21280 18991 21616 20021
rect 21280 18896 21372 18991
rect 21509 18896 21616 18991
rect 21280 17285 21616 18896
rect 21280 17212 21407 17285
rect 21487 17212 21616 17285
rect 21280 16191 21616 17212
rect 21280 16096 21381 16191
rect 21518 16096 21616 16191
rect 21280 14481 21616 16096
rect 21280 14410 21397 14481
rect 21484 14410 21616 14481
rect 21280 13390 21616 14410
rect 21280 13295 21385 13390
rect 21522 13295 21616 13390
rect 21280 11686 21616 13295
rect 21280 11610 21397 11686
rect 21483 11610 21616 11686
rect 21280 10586 21616 11610
rect 21280 10491 21370 10586
rect 21507 10491 21616 10586
rect 21280 8885 21616 10491
rect 21280 8811 21397 8885
rect 21484 8811 21616 8885
rect 21280 7791 21616 8811
rect 21280 7696 21374 7791
rect 21511 7696 21616 7791
rect 21280 6083 21616 7696
rect 21280 6011 21400 6083
rect 21485 6011 21616 6083
rect 21280 4985 21616 6011
rect 21280 4890 21381 4985
rect 21518 4890 21616 4985
rect 21280 3283 21616 4890
rect 21280 3212 21401 3283
rect 21486 3212 21616 3283
rect 21280 2186 21616 3212
rect 21280 2091 21382 2186
rect 21519 2091 21616 2186
rect 21280 480 21616 2091
rect 21280 408 21402 480
rect 21481 408 21616 480
rect 21280 198 21616 408
rect 16466 -327 16798 -252
rect 16466 -602 16535 -327
rect 16756 -602 16798 -327
rect 16466 -717 16798 -602
rect 18144 -1002 18483 123
rect 21279 56 21616 198
rect 23352 20944 23688 23184
rect 27776 23251 28112 27719
rect 27776 23179 27862 23251
rect 28000 23179 28112 23251
rect 23352 20862 23462 20944
rect 23576 20862 23688 20944
rect 23352 20151 23688 20862
rect 23352 20033 23421 20151
rect 23587 20033 23688 20151
rect 23352 18143 23688 20033
rect 23352 18068 23464 18143
rect 23575 18068 23688 18143
rect 23352 17275 23688 18068
rect 23352 17157 23416 17275
rect 23582 17157 23688 17275
rect 23352 15324 23688 17157
rect 23352 15258 23462 15324
rect 23577 15258 23688 15324
rect 23352 14424 23688 15258
rect 23352 14306 23431 14424
rect 23597 14306 23688 14424
rect 23352 12526 23688 14306
rect 23352 12460 23462 12526
rect 23577 12460 23688 12526
rect 23352 11689 23688 12460
rect 23352 11571 23442 11689
rect 23608 11571 23688 11689
rect 23352 9726 23688 11571
rect 23352 9663 23463 9726
rect 23578 9663 23688 9726
rect 23352 8900 23688 9663
rect 23352 8782 23446 8900
rect 23612 8782 23688 8900
rect 23352 6928 23688 8782
rect 23352 6865 23462 6928
rect 23577 6865 23688 6928
rect 23352 6175 23688 6865
rect 23352 6057 23435 6175
rect 23601 6057 23688 6175
rect 23352 4127 23688 6057
rect 23352 4056 23460 4127
rect 23576 4056 23688 4127
rect 23352 3330 23688 4056
rect 23352 3212 23433 3330
rect 23599 3212 23688 3330
rect 23352 2343 23688 3212
rect 26152 22456 26488 22632
rect 26152 22400 26292 22456
rect 26348 22400 26488 22456
rect 26152 21788 26488 22400
rect 26152 21693 26252 21788
rect 26389 21693 26488 21788
rect 26152 20089 26488 21693
rect 26152 20017 26277 20089
rect 26366 20017 26488 20089
rect 26152 18989 26488 20017
rect 26152 18894 26257 18989
rect 26394 18894 26488 18989
rect 26152 17285 26488 18894
rect 26152 17214 26270 17285
rect 26369 17214 26488 17285
rect 26152 16187 26488 17214
rect 26152 16092 26255 16187
rect 26392 16092 26488 16187
rect 26152 14483 26488 16092
rect 26152 14414 26265 14483
rect 26371 14414 26488 14483
rect 26152 13391 26488 14414
rect 26152 13296 26250 13391
rect 26387 13296 26488 13391
rect 26152 11687 26488 13296
rect 26152 11611 26278 11687
rect 26367 11611 26488 11687
rect 26152 10593 26488 11611
rect 26152 10498 26254 10593
rect 26391 10498 26488 10593
rect 26152 8886 26488 10498
rect 26152 8811 26265 8886
rect 26364 8811 26488 8886
rect 26152 7796 26488 8811
rect 26152 7701 26252 7796
rect 26389 7701 26488 7796
rect 26152 6090 26488 7701
rect 26152 6010 26275 6090
rect 26367 6010 26488 6090
rect 26152 4986 26488 6010
rect 26152 4891 26261 4986
rect 26398 4891 26488 4986
rect 26152 3290 26488 4891
rect 26152 3210 26264 3290
rect 26360 3210 26488 3290
rect 23352 1342 23690 2343
rect 23352 1271 23462 1342
rect 23578 1271 23690 1342
rect 23352 501 23690 1271
rect 23352 383 23406 501
rect 23572 383 23690 501
rect 21279 -252 21613 56
rect 23352 -252 23690 383
rect 21281 -414 21610 -252
rect 21281 -664 21332 -414
rect 21563 -664 21610 -414
rect 21281 -753 21610 -664
rect 23355 -1002 23690 -252
rect 26152 2188 26488 3210
rect 26152 2093 26252 2188
rect 26389 2093 26488 2188
rect 26152 483 26488 2093
rect 26152 406 26275 483
rect 26363 406 26488 483
rect 26152 180 26488 406
rect 27776 20937 28112 23179
rect 27776 20864 27887 20937
rect 28000 20864 28112 20937
rect 27776 20137 28112 20864
rect 27776 20019 27860 20137
rect 28026 20019 28112 20137
rect 27776 18139 28112 20019
rect 27776 18066 27889 18139
rect 28002 18066 28112 18139
rect 27776 17296 28112 18066
rect 27776 17178 27852 17296
rect 28018 17178 28112 17296
rect 27776 14428 28112 17178
rect 27776 14310 27862 14428
rect 28028 14310 28112 14428
rect 27776 12527 28112 14310
rect 27776 12456 27889 12527
rect 28001 12456 28112 12527
rect 27776 11712 28112 12456
rect 27776 11594 27865 11712
rect 28031 11594 28112 11712
rect 27776 9733 28112 11594
rect 27776 9663 27888 9733
rect 28000 9663 28112 9733
rect 27776 8887 28112 9663
rect 27776 8769 27859 8887
rect 28025 8769 28112 8887
rect 27776 6144 28112 8769
rect 27776 6026 27857 6144
rect 28023 6026 28112 6144
rect 27776 4123 28112 6026
rect 27776 4050 27887 4123
rect 28001 4050 28112 4123
rect 27776 3321 28112 4050
rect 27776 3203 27873 3321
rect 28039 3203 28112 3321
rect 27776 1330 28112 3203
rect 27776 1257 27887 1330
rect 28001 1257 28112 1330
rect 27776 474 28112 1257
rect 27776 356 27873 474
rect 28039 356 28112 474
rect 26152 -380 26491 180
rect 27776 -9 28112 356
rect 30968 22456 31304 22874
rect 30968 22400 31111 22456
rect 31167 22400 31304 22456
rect 30968 21793 31304 22400
rect 30968 21698 31071 21793
rect 31208 21698 31304 21793
rect 30968 20077 31304 21698
rect 30968 20020 31079 20077
rect 31192 20020 31304 20077
rect 30968 18990 31304 20020
rect 30968 18895 31066 18990
rect 31203 18895 31304 18990
rect 30968 17279 31304 18895
rect 30968 17221 31080 17279
rect 31192 17221 31304 17279
rect 30968 16191 31304 17221
rect 30968 16096 31065 16191
rect 31202 16096 31304 16191
rect 30968 14479 31304 16096
rect 30968 14423 31080 14479
rect 31192 14423 31304 14479
rect 30968 13393 31304 14423
rect 30968 13298 31068 13393
rect 31205 13298 31304 13393
rect 30968 11685 31304 13298
rect 30968 11625 31080 11685
rect 31192 11625 31304 11685
rect 30968 10594 31304 11625
rect 30968 10499 31064 10594
rect 31201 10499 31304 10594
rect 30968 8882 31304 10499
rect 30968 8826 31079 8882
rect 31192 8826 31304 8882
rect 30968 7792 31304 8826
rect 30968 7697 31063 7792
rect 31200 7697 31304 7792
rect 30968 6082 31304 7697
rect 30968 6026 31080 6082
rect 31193 6026 31304 6082
rect 30968 4994 31304 6026
rect 30968 4899 31065 4994
rect 31202 4899 31304 4994
rect 30968 3278 31304 4899
rect 30968 3222 31080 3278
rect 31192 3222 31304 3278
rect 30968 2197 31304 3222
rect 30968 2102 31069 2197
rect 31206 2102 31304 2197
rect 30968 482 31304 2102
rect 32928 20938 33264 27719
rect 32928 20874 33039 20938
rect 33155 20874 33264 20938
rect 32928 20146 33264 20874
rect 32928 20028 33016 20146
rect 33182 20028 33264 20146
rect 32928 18117 33264 20028
rect 32928 18053 33038 18117
rect 33154 18053 33264 18117
rect 32928 17287 33264 18053
rect 32928 17169 32994 17287
rect 33160 17169 33264 17287
rect 32928 15339 33264 17169
rect 32928 15269 33040 15339
rect 33152 15269 33264 15339
rect 32928 14433 33264 15269
rect 32928 14315 33000 14433
rect 33166 14315 33264 14433
rect 32928 12535 33264 14315
rect 32928 12465 33040 12535
rect 33152 12465 33264 12535
rect 32928 11686 33264 12465
rect 32928 11568 33008 11686
rect 33174 11568 33264 11686
rect 32928 9732 33264 11568
rect 32928 9666 33031 9732
rect 33143 9666 33264 9732
rect 32928 8891 33264 9666
rect 32928 8773 33001 8891
rect 33167 8773 33264 8891
rect 32928 6930 33264 8773
rect 32928 6864 33041 6930
rect 33153 6864 33264 6930
rect 32928 6141 33264 6864
rect 32928 6023 33030 6141
rect 33196 6023 33264 6141
rect 32928 4136 33264 6023
rect 32928 4072 33030 4136
rect 33139 4072 33264 4136
rect 32928 3332 33264 4072
rect 32928 3214 33004 3332
rect 33170 3214 33264 3332
rect 32928 1329 33264 3214
rect 32928 1265 33043 1329
rect 33152 1265 33264 1329
rect 35672 26199 36008 27719
rect 35672 26137 35783 26199
rect 35896 26137 36008 26199
rect 35672 25238 36008 26137
rect 35672 25176 35784 25238
rect 35897 25176 36008 25238
rect 35672 24283 36008 25176
rect 35672 24221 35784 24283
rect 35896 24221 36008 24283
rect 35672 23300 36008 24221
rect 35672 23238 35784 23300
rect 35896 23238 36008 23300
rect 35672 20928 36008 23238
rect 35672 20869 35784 20928
rect 35896 20869 36008 20928
rect 35672 20145 36008 20869
rect 35672 20027 35763 20145
rect 35929 20027 36008 20145
rect 35672 18127 36008 20027
rect 35672 18068 35784 18127
rect 35896 18068 36008 18127
rect 35672 17298 36008 18068
rect 35672 17180 35768 17298
rect 35934 17180 36008 17298
rect 35672 15333 36008 17180
rect 35672 15274 35784 15333
rect 35896 15274 36008 15333
rect 35672 14446 36008 15274
rect 35672 14328 35761 14446
rect 35927 14328 36008 14446
rect 35672 12524 36008 14328
rect 35672 12465 35784 12524
rect 35896 12465 36008 12524
rect 35672 11693 36008 12465
rect 35672 11575 35764 11693
rect 35930 11575 36008 11693
rect 35672 9732 36008 11575
rect 35672 9674 35784 9732
rect 35896 9674 36008 9732
rect 35672 8896 36008 9674
rect 35672 8778 35758 8896
rect 35924 8778 36008 8896
rect 35672 6921 36008 8778
rect 35672 6863 35784 6921
rect 35896 6863 36008 6921
rect 35672 6142 36008 6863
rect 35672 6024 35754 6142
rect 35920 6024 36008 6142
rect 35672 4130 36008 6024
rect 35672 4074 35783 4130
rect 35896 4074 36008 4130
rect 35672 3368 36008 4074
rect 35672 3250 35753 3368
rect 35919 3250 36008 3368
rect 35672 1322 36008 3250
rect 32928 740 33264 1265
rect 30968 421 31079 482
rect 31193 421 31304 482
rect 30968 74 31304 421
rect 27776 -224 28113 -9
rect 26152 -637 26205 -380
rect 26428 -637 26491 -380
rect 26152 -704 26491 -637
rect 27778 -1002 28113 -224
rect 30967 -112 31304 74
rect 32921 492 33264 740
rect 32921 374 33018 492
rect 33184 374 33264 492
rect 32921 -56 33264 374
rect 35671 492 36008 1322
rect 35671 374 35762 492
rect 35928 374 36008 492
rect 35671 -56 36008 374
rect 37016 25450 37352 26600
rect 37016 25297 37069 25450
rect 37310 25297 37352 25450
rect 37016 24500 37352 25297
rect 37016 24347 37073 24500
rect 37314 24347 37352 24500
rect 37016 23532 37352 24347
rect 37016 23379 37061 23532
rect 37302 23379 37352 23532
rect 37016 22563 37352 23379
rect 37016 22410 37071 22563
rect 37312 22410 37352 22563
rect 37016 21790 37352 22410
rect 37016 21695 37117 21790
rect 37254 21695 37352 21790
rect 37016 20089 37352 21695
rect 37016 20023 37145 20089
rect 37223 20023 37352 20089
rect 37016 18993 37352 20023
rect 37016 18898 37124 18993
rect 37261 18898 37352 18993
rect 37016 17289 37352 18898
rect 37016 17220 37143 17289
rect 37219 17220 37352 17289
rect 37016 16191 37352 17220
rect 37016 16096 37119 16191
rect 37256 16096 37352 16191
rect 37016 14489 37352 16096
rect 37016 14425 37150 14489
rect 37224 14425 37352 14489
rect 37016 13391 37352 14425
rect 37016 13296 37119 13391
rect 37256 13296 37352 13391
rect 37016 11686 37352 13296
rect 37016 11618 37146 11686
rect 37224 11618 37352 11686
rect 37016 10590 37352 11618
rect 37016 10495 37110 10590
rect 37247 10495 37352 10590
rect 37016 8885 37352 10495
rect 37016 8812 37142 8885
rect 37224 8812 37352 8885
rect 37016 7792 37352 8812
rect 37016 7697 37118 7792
rect 37255 7697 37352 7792
rect 37016 6083 37352 7697
rect 37016 6015 37140 6083
rect 37224 6015 37352 6083
rect 37016 4990 37352 6015
rect 37016 4895 37116 4990
rect 37253 4895 37352 4990
rect 37016 3285 37352 4895
rect 37016 3219 37137 3285
rect 37225 3219 37352 3285
rect 37016 2151 37352 3219
rect 44397 20330 46986 27719
rect 44397 19881 45369 20330
rect 46227 19881 46986 20330
rect 44397 17465 46986 19881
rect 44397 17026 45342 17465
rect 46161 17026 46986 17465
rect 44397 14587 46986 17026
rect 44397 14190 45345 14587
rect 46149 14190 46986 14587
rect 44397 11854 46986 14190
rect 44397 11435 45276 11854
rect 46096 11435 46986 11854
rect 44397 9063 46986 11435
rect 44397 8662 45317 9063
rect 46126 8662 46986 9063
rect 44397 6288 46986 8662
rect 44397 5920 45246 6288
rect 46070 5920 46986 6288
rect 44397 3499 46986 5920
rect 44397 3119 45192 3499
rect 46104 3119 46986 3499
rect 44397 2362 46986 3119
rect 37016 2056 37117 2151
rect 37254 2056 37352 2151
rect 37016 -56 37352 2056
rect 30967 -252 31301 -112
rect 30967 -393 31300 -252
rect 30967 -662 31011 -393
rect 31255 -662 31300 -393
rect 30967 -754 31300 -662
rect -2581 -1006 28113 -1002
rect 32921 -1006 33262 -56
rect 35671 -1006 36007 -56
rect 37018 -252 37352 -56
rect 44397 663 46986 1899
rect 44397 245 45293 663
rect 46226 245 46986 663
rect 37019 -368 37350 -252
rect 44397 -259 46986 245
rect 37019 -659 37051 -368
rect 37326 -659 37350 -368
rect 37019 -775 37350 -659
rect 44390 -1006 46988 -259
rect -2581 -1009 46988 -1006
rect -6204 -3591 46988 -1009
rect -6204 -3592 -312 -3591
rect 27800 -3594 46988 -3591
rect 44390 -3597 46988 -3594
<< via4 >>
rect -5232 20293 -4434 20317
rect -5297 19920 -4423 20293
rect -5232 19913 -4434 19920
rect -5228 17031 -4377 17438
rect -5317 14179 -4466 14586
rect -5253 11443 -4402 11850
rect -5326 8639 -4475 9046
rect -5235 5902 -4384 6309
rect -5349 3098 -4498 3505
rect 364 20027 530 20145
rect 359 17180 525 17298
rect 362 14310 528 14428
rect 365 11591 531 11709
rect 369 8783 535 8901
rect 370 6033 536 6151
rect 364 3234 530 3352
rect 2169 21777 2306 21788
rect 2169 21703 2184 21777
rect 2184 21703 2296 21777
rect 2296 21703 2306 21777
rect 2169 21693 2306 21703
rect 2169 18973 2306 18988
rect 2169 18907 2184 18973
rect 2184 18907 2296 18973
rect 2296 18907 2306 18973
rect 2169 18893 2306 18907
rect 2171 16181 2308 16197
rect 2171 16117 2184 16181
rect 2184 16117 2296 16181
rect 2296 16117 2308 16181
rect 2171 16102 2308 16117
rect 2175 13383 2312 13393
rect 2175 13310 2184 13383
rect 2184 13310 2296 13383
rect 2296 13310 2312 13383
rect 2175 13298 2312 13310
rect 2172 10581 2309 10591
rect 2172 10503 2184 10581
rect 2184 10503 2296 10581
rect 2296 10503 2309 10581
rect 2172 10496 2309 10503
rect 2170 7784 2307 7795
rect 2170 7714 2184 7784
rect 2184 7714 2296 7784
rect 2296 7714 2307 7784
rect 2170 7700 2307 7714
rect 2173 4984 2310 4995
rect 2173 4910 2184 4984
rect 2184 4910 2296 4984
rect 2296 4910 2310 4984
rect 2173 4900 2310 4910
rect 2171 2172 2308 2187
rect 2171 2104 2184 2172
rect 2184 2104 2296 2172
rect 2296 2104 2308 2172
rect 2171 2092 2308 2104
rect -5047 246 -4196 653
rect 359 371 525 489
rect 3835 20021 4001 20139
rect 3826 17164 3992 17282
rect 3830 14323 3996 14441
rect 3841 11590 4007 11708
rect 3834 8769 4000 8887
rect 3825 6023 3991 6141
rect 3837 3221 4003 3339
rect 3831 384 3997 502
rect 6877 21776 7014 21787
rect 6877 21698 6887 21776
rect 6887 21698 7001 21776
rect 7001 21698 7014 21776
rect 6877 21692 7014 21698
rect 6875 18976 7012 18988
rect 6875 18901 6888 18976
rect 6888 18901 7000 18976
rect 7000 18901 7012 18976
rect 6875 18893 7012 18901
rect 6873 16173 7010 16186
rect 6873 16104 6887 16173
rect 6887 16104 7000 16173
rect 7000 16104 7010 16173
rect 6873 16091 7010 16104
rect 6871 13374 7008 13388
rect 6871 13305 6885 13374
rect 6885 13305 7001 13374
rect 7001 13305 7008 13374
rect 6871 13293 7008 13305
rect 6876 10576 7013 10592
rect 6876 10505 6887 10576
rect 6887 10505 7001 10576
rect 7001 10505 7013 10576
rect 6876 10497 7013 10505
rect 6872 7773 7009 7787
rect 6872 7708 6888 7773
rect 6888 7708 7000 7773
rect 7000 7708 7009 7773
rect 6872 7692 7009 7708
rect 6872 4974 7009 4990
rect 6872 4903 6888 4974
rect 6888 4903 7001 4974
rect 7001 4903 7009 4974
rect 6872 4895 7009 4903
rect 6874 2173 7011 2190
rect 6874 2104 6887 2173
rect 6887 2104 7001 2173
rect 7001 2104 7011 2173
rect 6874 2095 7011 2104
rect 2128 -657 2367 -402
rect 8650 20043 8816 20161
rect 8652 17166 8818 17284
rect 8642 14319 8808 14437
rect 8663 11578 8829 11696
rect 8649 8769 8815 8887
rect 8664 6019 8830 6137
rect 8657 3239 8823 3357
rect 8648 365 8814 483
rect 11750 21782 11887 21791
rect 11750 21700 11760 21782
rect 11760 21700 11873 21782
rect 11873 21700 11887 21782
rect 11750 21696 11887 21700
rect 11745 18986 11882 18989
rect 11745 18904 11760 18986
rect 11760 18904 11872 18986
rect 11872 18904 11882 18986
rect 11745 18894 11882 18904
rect 11748 16180 11885 16192
rect 11748 16110 11762 16180
rect 11762 16110 11873 16180
rect 11873 16110 11885 16180
rect 11748 16097 11885 16110
rect 11743 13384 11880 13394
rect 11743 13308 11760 13384
rect 11760 13308 11873 13384
rect 11873 13308 11880 13384
rect 11743 13299 11880 13308
rect 11745 10583 11882 10589
rect 11745 10508 11760 10583
rect 11760 10508 11872 10583
rect 11872 10508 11882 10583
rect 11745 10494 11882 10508
rect 11746 7781 11883 7789
rect 11746 7703 11760 7781
rect 11760 7703 11872 7781
rect 11872 7703 11883 7781
rect 11746 7694 11883 7703
rect 11745 4980 11882 4991
rect 11745 4907 11759 4980
rect 11759 4907 11872 4980
rect 11872 4907 11882 4980
rect 11745 4896 11882 4907
rect 13853 20019 14019 20137
rect 13849 17175 14015 17293
rect 13851 14308 14017 14426
rect 13858 11605 14024 11723
rect 13869 8773 14035 8891
rect 13856 6014 14022 6132
rect 13858 3236 14024 3354
rect 16568 21769 16705 21791
rect 16568 21710 16593 21769
rect 16593 21710 16683 21769
rect 16683 21710 16705 21769
rect 16568 21696 16705 21710
rect 16563 18969 16700 18989
rect 16563 18910 16593 18969
rect 16593 18910 16665 18969
rect 16665 18910 16700 18969
rect 16563 18894 16700 18910
rect 16561 16175 16698 16194
rect 16561 16114 16588 16175
rect 16588 16114 16667 16175
rect 16667 16114 16698 16175
rect 16561 16099 16698 16114
rect 16562 13372 16699 13393
rect 16562 13308 16594 13372
rect 16594 13308 16668 13372
rect 16668 13308 16699 13372
rect 16562 13298 16699 13308
rect 16565 10574 16702 10594
rect 16565 10512 16593 10574
rect 16593 10512 16669 10574
rect 16669 10512 16702 10574
rect 16565 10499 16702 10512
rect 16561 7772 16698 7790
rect 16561 7706 16589 7772
rect 16589 7706 16670 7772
rect 16670 7706 16698 7772
rect 16561 7695 16698 7706
rect 16561 4976 16698 4984
rect 16561 4906 16589 4976
rect 16589 4906 16672 4976
rect 16672 4906 16698 4976
rect 16561 4889 16698 4906
rect 11748 2181 11885 2191
rect 11748 2106 11758 2181
rect 11758 2106 11876 2181
rect 11876 2106 11885 2181
rect 11748 2096 11885 2106
rect 6823 -696 7082 -431
rect 13863 366 14029 484
rect 11709 -606 11938 -393
rect 16565 2177 16702 2190
rect 16565 2104 16595 2177
rect 16595 2104 16675 2177
rect 16675 2104 16702 2177
rect 16565 2095 16702 2104
rect 18229 20024 18395 20142
rect 18202 17157 18368 17275
rect 18237 14315 18403 14433
rect 18236 11571 18402 11689
rect 18240 8773 18406 8891
rect 18232 6028 18398 6146
rect 18226 3240 18392 3358
rect 18221 381 18387 499
rect 21386 21773 21523 21788
rect 21386 21709 21412 21773
rect 21412 21709 21490 21773
rect 21490 21709 21523 21773
rect 21386 21693 21523 21709
rect 21372 18978 21509 18991
rect 21372 18914 21404 18978
rect 21404 18914 21481 18978
rect 21481 18914 21509 18978
rect 21372 18896 21509 18914
rect 21381 16181 21518 16191
rect 21381 16108 21411 16181
rect 21411 16108 21491 16181
rect 21491 16108 21518 16181
rect 21381 16096 21518 16108
rect 21385 13376 21522 13390
rect 21385 13305 21406 13376
rect 21406 13305 21493 13376
rect 21493 13305 21522 13376
rect 21385 13295 21522 13305
rect 21370 10576 21507 10586
rect 21370 10500 21402 10576
rect 21402 10500 21488 10576
rect 21488 10500 21507 10576
rect 21370 10491 21507 10500
rect 21374 7779 21511 7791
rect 21374 7705 21404 7779
rect 21404 7705 21491 7779
rect 21491 7705 21511 7779
rect 21374 7696 21511 7705
rect 21381 4974 21518 4985
rect 21381 4902 21408 4974
rect 21408 4902 21493 4974
rect 21493 4902 21518 4974
rect 21381 4890 21518 4902
rect 21382 2174 21519 2186
rect 21382 2103 21403 2174
rect 21403 2103 21488 2174
rect 21488 2103 21519 2174
rect 21382 2091 21519 2103
rect 16535 -602 16756 -327
rect 23421 20033 23587 20151
rect 23416 17157 23582 17275
rect 23431 14306 23597 14424
rect 23442 11571 23608 11689
rect 23446 8782 23612 8900
rect 23435 6057 23601 6175
rect 23433 3212 23599 3330
rect 26252 21776 26389 21788
rect 26252 21706 26264 21776
rect 26264 21706 26375 21776
rect 26375 21706 26389 21776
rect 26252 21693 26389 21706
rect 26257 18975 26394 18989
rect 26257 18903 26281 18975
rect 26281 18903 26370 18975
rect 26370 18903 26394 18975
rect 26257 18894 26394 18903
rect 26255 16176 26392 16187
rect 26255 16105 26271 16176
rect 26271 16105 26370 16176
rect 26370 16105 26392 16176
rect 26255 16092 26392 16105
rect 26250 13380 26387 13391
rect 26250 13311 26267 13380
rect 26267 13311 26373 13380
rect 26373 13311 26387 13380
rect 26250 13296 26387 13311
rect 26254 10582 26391 10593
rect 26254 10506 26277 10582
rect 26277 10506 26366 10582
rect 26366 10506 26391 10582
rect 26254 10498 26391 10506
rect 26252 7783 26389 7796
rect 26252 7708 26273 7783
rect 26273 7708 26372 7783
rect 26372 7708 26389 7783
rect 26252 7701 26389 7708
rect 26261 4980 26398 4986
rect 26261 4900 26281 4980
rect 26281 4900 26373 4980
rect 26373 4900 26398 4980
rect 26261 4891 26398 4900
rect 23406 383 23572 501
rect 21332 -664 21563 -414
rect 26252 2179 26389 2188
rect 26252 2099 26276 2179
rect 26276 2099 26372 2179
rect 26372 2099 26389 2179
rect 26252 2093 26389 2099
rect 27860 20019 28026 20137
rect 27852 17178 28018 17296
rect 27862 14310 28028 14428
rect 27865 11594 28031 11712
rect 27859 8769 28025 8887
rect 27857 6026 28023 6144
rect 27873 3203 28039 3321
rect 27873 356 28039 474
rect 31071 21771 31208 21793
rect 31071 21714 31080 21771
rect 31080 21714 31193 21771
rect 31193 21714 31208 21771
rect 31071 21698 31208 21714
rect 31066 18969 31203 18990
rect 31066 18911 31080 18969
rect 31080 18911 31192 18969
rect 31192 18911 31203 18969
rect 31066 18895 31203 18911
rect 31065 16171 31202 16191
rect 31065 16115 31080 16171
rect 31080 16115 31192 16171
rect 31192 16115 31202 16171
rect 31065 16096 31202 16115
rect 31068 13370 31205 13393
rect 31068 13310 31080 13370
rect 31080 13310 31192 13370
rect 31192 13310 31205 13370
rect 31068 13298 31205 13310
rect 31064 10574 31201 10594
rect 31064 10518 31080 10574
rect 31080 10518 31193 10574
rect 31193 10518 31201 10574
rect 31064 10499 31201 10518
rect 31063 7772 31200 7792
rect 31063 7716 31079 7772
rect 31079 7716 31192 7772
rect 31192 7716 31200 7772
rect 31063 7697 31200 7716
rect 31065 4977 31202 4994
rect 31065 4921 31080 4977
rect 31080 4921 31192 4977
rect 31192 4921 31202 4977
rect 31065 4899 31202 4921
rect 31069 2178 31206 2197
rect 31069 2117 31079 2178
rect 31079 2117 31193 2178
rect 31193 2117 31206 2178
rect 31069 2102 31206 2117
rect 33016 20028 33182 20146
rect 32994 17169 33160 17287
rect 33000 14315 33166 14433
rect 33008 11568 33174 11686
rect 33001 8773 33167 8891
rect 33030 6023 33196 6141
rect 33004 3214 33170 3332
rect 35763 20027 35929 20145
rect 35768 17180 35934 17298
rect 35761 14328 35927 14446
rect 35764 11575 35930 11693
rect 35758 8778 35924 8896
rect 35754 6024 35920 6142
rect 35753 3250 35919 3368
rect 26205 -637 26428 -380
rect 33018 374 33184 492
rect 35762 374 35928 492
rect 37069 25411 37310 25450
rect 37069 25335 37139 25411
rect 37139 25335 37230 25411
rect 37230 25335 37310 25411
rect 37069 25297 37310 25335
rect 37073 24454 37314 24500
rect 37073 24378 37137 24454
rect 37137 24378 37228 24454
rect 37228 24378 37314 24454
rect 37073 24347 37314 24378
rect 37061 23495 37302 23532
rect 37061 23426 37140 23495
rect 37140 23426 37220 23495
rect 37220 23426 37302 23495
rect 37061 23379 37302 23426
rect 37071 22518 37312 22563
rect 37071 22449 37137 22518
rect 37137 22449 37217 22518
rect 37217 22449 37312 22518
rect 37071 22410 37312 22449
rect 37117 21773 37254 21790
rect 37117 21707 37146 21773
rect 37146 21707 37224 21773
rect 37224 21707 37254 21773
rect 37117 21695 37254 21707
rect 37124 18978 37261 18993
rect 37124 18909 37151 18978
rect 37151 18909 37227 18978
rect 37227 18909 37261 18978
rect 37124 18898 37261 18909
rect 37119 16175 37256 16191
rect 37119 16111 37144 16175
rect 37144 16111 37218 16175
rect 37218 16111 37256 16175
rect 37119 16096 37256 16111
rect 37119 13376 37256 13391
rect 37119 13308 37148 13376
rect 37148 13308 37226 13376
rect 37226 13308 37256 13376
rect 37119 13296 37256 13308
rect 37110 10579 37247 10590
rect 37110 10506 37137 10579
rect 37137 10506 37219 10579
rect 37219 10506 37247 10579
rect 37110 10495 37247 10506
rect 37118 7779 37255 7792
rect 37118 7711 37144 7779
rect 37144 7711 37228 7779
rect 37228 7711 37255 7779
rect 37118 7697 37255 7711
rect 37116 4976 37253 4990
rect 37116 4910 37140 4976
rect 37140 4910 37228 4976
rect 37228 4910 37253 4976
rect 37116 4895 37253 4910
rect 45369 19881 46227 20330
rect 45342 17026 46161 17465
rect 45345 14190 46149 14587
rect 45276 11435 46096 11854
rect 45317 8662 46126 9063
rect 45246 5920 46070 6288
rect 45192 3119 46104 3499
rect 37117 2056 37254 2151
rect 31011 -662 31255 -393
rect 45293 245 46226 663
rect 37051 -659 37326 -368
<< metal5 >>
rect 16466 34813 16800 34815
rect -7281 34812 21156 34813
rect 22595 34812 26507 34813
rect -7281 34810 51435 34812
rect -9848 32224 51435 34810
rect -9848 28871 -7264 32224
rect -9849 22018 -7261 28871
rect -9849 22007 -1615 22018
rect 2073 22007 2408 32224
rect -9849 22004 6503 22007
rect 6777 22004 7111 32224
rect 11648 24623 11982 32224
rect 11648 22996 11981 24623
rect 16466 24611 16800 32224
rect 11648 22007 11982 22996
rect 16466 22700 16798 24611
rect 16466 22007 16800 22700
rect 21282 22007 21614 32224
rect 26154 32223 51435 32224
rect 26154 22007 26486 32223
rect 30968 22007 31300 32223
rect 37017 25450 37349 32223
rect 37017 25297 37069 25450
rect 37310 25297 37349 25450
rect 37017 24500 37349 25297
rect 37017 24347 37073 24500
rect 37314 24347 37349 24500
rect 37017 23532 37349 24347
rect 37017 23379 37061 23532
rect 37302 23379 37349 23532
rect 37017 22563 37349 23379
rect 37017 22410 37071 22563
rect 37312 22410 37349 22563
rect 37017 22007 37349 22410
rect 48849 31739 51435 32223
rect 48849 29599 51437 31739
rect 48849 22019 51439 29599
rect 42427 22007 51439 22019
rect 7343 22004 51439 22007
rect -9849 21793 51439 22004
rect -9849 21791 31071 21793
rect -9849 21788 11750 21791
rect -9849 21693 2169 21788
rect 2306 21787 11750 21788
rect 2306 21693 6877 21787
rect -9849 21692 6877 21693
rect 7014 21696 11750 21787
rect 11887 21696 16568 21791
rect 16705 21788 31071 21791
rect 16705 21696 21386 21788
rect 7014 21693 21386 21696
rect 21523 21693 26252 21788
rect 26389 21698 31071 21788
rect 31208 21790 51439 21793
rect 31208 21698 37117 21790
rect 26389 21695 37117 21698
rect 37254 21695 51439 21790
rect 26389 21693 51439 21695
rect 7014 21692 51439 21693
rect -9849 21560 51439 21692
rect -9849 21555 -1615 21560
rect 42427 21556 51439 21560
rect -9849 19163 -7261 21555
rect -5616 20327 -1762 20332
rect 43111 20330 46517 20332
rect 43111 20328 45369 20330
rect 42896 20327 45369 20328
rect -5616 20317 45369 20327
rect -5616 20293 -5232 20317
rect -4434 20293 45369 20317
rect -5616 19920 -5297 20293
rect -4423 20161 45369 20293
rect -4423 20145 8650 20161
rect -4423 20027 364 20145
rect 530 20139 8650 20145
rect 530 20027 3835 20139
rect -4423 20021 3835 20027
rect 4001 20043 8650 20139
rect 8816 20151 45369 20161
rect 8816 20142 23421 20151
rect 8816 20137 18229 20142
rect 8816 20043 13853 20137
rect 4001 20021 13853 20043
rect -4423 20019 13853 20021
rect 14019 20024 18229 20137
rect 18395 20033 23421 20142
rect 23587 20146 45369 20151
rect 23587 20137 33016 20146
rect 23587 20033 27860 20137
rect 18395 20024 27860 20033
rect 14019 20019 27860 20024
rect 28026 20028 33016 20137
rect 33182 20145 45369 20146
rect 33182 20028 35763 20145
rect 28026 20027 35763 20028
rect 35929 20027 45369 20145
rect 28026 20019 45369 20027
rect -4423 19920 45369 20019
rect -5616 19913 -5232 19920
rect -4434 19913 45369 19920
rect -5616 19881 45369 19913
rect 46227 19881 46517 20330
rect -5616 19880 46517 19881
rect -5616 19879 -1762 19880
rect -9849 19151 -1259 19163
rect 48849 19161 51439 21556
rect 42557 19151 51439 19161
rect -9849 18993 51439 19151
rect -9849 18991 37124 18993
rect -9849 18989 21372 18991
rect -9849 18988 11745 18989
rect -9849 18893 2169 18988
rect 2306 18893 6875 18988
rect 7012 18894 11745 18988
rect 11882 18894 16563 18989
rect 16700 18896 21372 18989
rect 21509 18990 37124 18991
rect 21509 18989 31066 18990
rect 21509 18896 26257 18989
rect 16700 18894 26257 18896
rect 26394 18895 31066 18989
rect 31203 18898 37124 18990
rect 37261 18898 51439 18993
rect 31203 18895 51439 18898
rect 26394 18894 51439 18895
rect 7012 18893 51439 18894
rect -9849 18704 51439 18893
rect -9849 18700 -1259 18704
rect -9849 16413 -7261 18700
rect 42557 18698 51439 18704
rect -5657 17471 -1803 17474
rect 42776 17471 43159 17472
rect -5657 17465 46877 17471
rect -5657 17438 45342 17465
rect -5657 17031 -5228 17438
rect -4377 17298 45342 17438
rect -4377 17180 359 17298
rect 525 17296 35768 17298
rect 525 17293 27852 17296
rect 525 17284 13849 17293
rect 525 17282 8652 17284
rect 525 17180 3826 17282
rect -4377 17164 3826 17180
rect 3992 17166 8652 17282
rect 8818 17175 13849 17284
rect 14015 17275 27852 17293
rect 14015 17175 18202 17275
rect 8818 17166 18202 17175
rect 3992 17164 18202 17166
rect -4377 17157 18202 17164
rect 18368 17157 23416 17275
rect 23582 17178 27852 17275
rect 28018 17287 35768 17296
rect 28018 17178 32994 17287
rect 23582 17169 32994 17178
rect 33160 17180 35768 17287
rect 35934 17180 45342 17298
rect 33160 17169 45342 17180
rect 23582 17157 45342 17169
rect -4377 17031 45342 17157
rect -5657 17026 45342 17031
rect 46161 17026 46877 17465
rect -5657 17024 46877 17026
rect -5657 17021 -1803 17024
rect 42986 17023 46877 17024
rect 48849 16429 51439 18698
rect -9849 16407 -1693 16413
rect 42733 16407 51439 16429
rect -9849 16197 51439 16407
rect -9849 16102 2171 16197
rect 2308 16194 51439 16197
rect 2308 16192 16561 16194
rect 2308 16186 11748 16192
rect 2308 16102 6873 16186
rect -9849 16091 6873 16102
rect 7010 16097 11748 16186
rect 11885 16099 16561 16192
rect 16698 16191 51439 16194
rect 16698 16099 21381 16191
rect 11885 16097 21381 16099
rect 7010 16096 21381 16097
rect 21518 16187 31065 16191
rect 21518 16096 26255 16187
rect 7010 16092 26255 16096
rect 26392 16096 31065 16187
rect 31202 16096 37119 16191
rect 37256 16096 51439 16191
rect 26392 16092 51439 16096
rect 7010 16091 51439 16092
rect -9849 15966 51439 16091
rect -9849 15960 42898 15966
rect -9849 15950 -1693 15960
rect -9849 13553 -7261 15950
rect -5701 14615 -1847 14619
rect 42990 14616 46591 14617
rect 42786 14615 46591 14616
rect -5701 14587 46591 14615
rect -5701 14586 45345 14587
rect -5701 14179 -5317 14586
rect -4466 14446 45345 14586
rect -4466 14441 35761 14446
rect -4466 14428 3830 14441
rect -4466 14310 362 14428
rect 528 14323 3830 14428
rect 3996 14437 35761 14441
rect 3996 14323 8642 14437
rect 528 14319 8642 14323
rect 8808 14433 35761 14437
rect 8808 14426 18237 14433
rect 8808 14319 13851 14426
rect 528 14310 13851 14319
rect -4466 14308 13851 14310
rect 14017 14315 18237 14426
rect 18403 14428 33000 14433
rect 18403 14424 27862 14428
rect 18403 14315 23431 14424
rect 14017 14308 23431 14315
rect -4466 14306 23431 14308
rect 23597 14310 27862 14424
rect 28028 14315 33000 14428
rect 33166 14328 35761 14433
rect 35927 14328 45345 14446
rect 33166 14315 45345 14328
rect 28028 14310 45345 14315
rect 23597 14306 45345 14310
rect -4466 14190 45345 14306
rect 46149 14190 46591 14587
rect -4466 14179 46591 14190
rect -5701 14168 46591 14179
rect -5701 14166 -1847 14168
rect 42990 14166 46591 14168
rect 48849 13567 51439 15966
rect -9849 13551 -1737 13553
rect 42753 13551 51439 13567
rect -9849 13394 51439 13551
rect -9849 13393 11743 13394
rect -9849 13298 2175 13393
rect 2312 13388 11743 13393
rect 2312 13298 6871 13388
rect -9849 13293 6871 13298
rect 7008 13299 11743 13388
rect 11880 13393 51439 13394
rect 11880 13299 16562 13393
rect 7008 13298 16562 13299
rect 16699 13391 31068 13393
rect 16699 13390 26250 13391
rect 16699 13298 21385 13390
rect 7008 13295 21385 13298
rect 21522 13296 26250 13390
rect 26387 13298 31068 13391
rect 31205 13391 51439 13393
rect 31205 13298 37119 13391
rect 26387 13296 37119 13298
rect 37256 13296 51439 13391
rect 21522 13295 51439 13296
rect 7008 13293 51439 13295
rect -9849 13104 51439 13293
rect -9849 13090 -1737 13104
rect -9849 10698 -7261 13090
rect -5588 11871 -1734 11873
rect 42661 11871 46558 11874
rect -5588 11854 46558 11871
rect -5588 11850 45276 11854
rect -5588 11443 -5253 11850
rect -4402 11723 45276 11850
rect -4402 11709 13858 11723
rect -4402 11591 365 11709
rect 531 11708 13858 11709
rect 531 11591 3841 11708
rect -4402 11590 3841 11591
rect 4007 11696 13858 11708
rect 4007 11590 8663 11696
rect -4402 11578 8663 11590
rect 8829 11605 13858 11696
rect 14024 11712 45276 11723
rect 14024 11689 27865 11712
rect 14024 11605 18236 11689
rect 8829 11578 18236 11605
rect -4402 11571 18236 11578
rect 18402 11571 23442 11689
rect 23608 11594 27865 11689
rect 28031 11693 45276 11712
rect 28031 11686 35764 11693
rect 28031 11594 33008 11686
rect 23608 11571 33008 11594
rect -4402 11568 33008 11571
rect 33174 11575 35764 11686
rect 35930 11575 45276 11693
rect 33174 11568 45276 11575
rect -4402 11443 45276 11568
rect -5588 11435 45276 11443
rect 46096 11435 46558 11854
rect -5588 11424 46558 11435
rect -5588 11420 -1734 11424
rect 42661 11419 46558 11424
rect 48849 10715 51439 13104
rect -9849 10695 -1778 10698
rect 42658 10695 51439 10715
rect -9849 10594 51439 10695
rect -9849 10592 16565 10594
rect -9849 10591 6876 10592
rect -9849 10496 2172 10591
rect 2309 10497 6876 10591
rect 7013 10589 16565 10592
rect 7013 10497 11745 10589
rect 2309 10496 11745 10497
rect -9849 10494 11745 10496
rect 11882 10499 16565 10589
rect 16702 10593 31064 10594
rect 16702 10586 26254 10593
rect 16702 10499 21370 10586
rect 11882 10494 21370 10499
rect -9849 10491 21370 10494
rect 21507 10498 26254 10586
rect 26391 10499 31064 10593
rect 31201 10590 51439 10594
rect 31201 10499 37110 10590
rect 26391 10498 37110 10499
rect 21507 10495 37110 10498
rect 37247 10495 51439 10590
rect 21507 10491 51439 10495
rect -9849 10252 51439 10491
rect -9849 10248 42898 10252
rect -9849 10235 -1778 10248
rect -9849 7958 -7261 10235
rect 42827 9071 46546 9074
rect -2352 9068 46546 9071
rect -5697 9063 46546 9068
rect -5697 9046 45317 9063
rect -5697 8639 -5326 9046
rect -4475 8901 45317 9046
rect -4475 8783 369 8901
rect 535 8900 45317 8901
rect 535 8891 23446 8900
rect 535 8887 13869 8891
rect 535 8783 3834 8887
rect -4475 8769 3834 8783
rect 4000 8769 8649 8887
rect 8815 8773 13869 8887
rect 14035 8773 18240 8891
rect 18406 8782 23446 8891
rect 23612 8896 45317 8900
rect 23612 8891 35758 8896
rect 23612 8887 33001 8891
rect 23612 8782 27859 8887
rect 18406 8773 27859 8782
rect 8815 8769 27859 8773
rect 28025 8773 33001 8887
rect 33167 8778 35758 8891
rect 35924 8778 45317 8896
rect 33167 8773 45317 8778
rect 28025 8769 45317 8773
rect -4475 8662 45317 8769
rect 46126 8662 46546 9063
rect -4475 8639 46546 8662
rect -5697 8625 46546 8639
rect -5697 8624 43159 8625
rect -5697 8623 -1806 8624
rect 42861 8622 43159 8624
rect 48849 7970 51439 10252
rect -9849 7951 -1866 7958
rect 42720 7951 51439 7970
rect -9849 7796 51439 7951
rect -9849 7795 26252 7796
rect -9849 7700 2170 7795
rect 2307 7791 26252 7795
rect 2307 7790 21374 7791
rect 2307 7789 16561 7790
rect 2307 7787 11746 7789
rect 2307 7700 6872 7787
rect -9849 7692 6872 7700
rect 7009 7694 11746 7787
rect 11883 7695 16561 7789
rect 16698 7696 21374 7790
rect 21511 7701 26252 7791
rect 26389 7792 51439 7796
rect 26389 7701 31063 7792
rect 21511 7697 31063 7701
rect 31200 7697 37118 7792
rect 37255 7697 51439 7792
rect 21511 7696 51439 7697
rect 16698 7695 51439 7696
rect 11883 7694 51439 7695
rect 7009 7692 51439 7694
rect -9849 7507 51439 7692
rect -9849 7504 42896 7507
rect -9849 7495 -1866 7504
rect -9849 5224 -7261 7495
rect 42823 6329 45612 6330
rect 42823 6327 46513 6329
rect -2352 6325 46513 6327
rect -5587 6309 46513 6325
rect -5587 5902 -5235 6309
rect -4384 6288 46513 6309
rect -4384 6175 45246 6288
rect -4384 6151 23435 6175
rect -4384 6033 370 6151
rect 536 6146 23435 6151
rect 536 6141 18232 6146
rect 536 6033 3825 6141
rect -4384 6023 3825 6033
rect 3991 6137 18232 6141
rect 3991 6023 8664 6137
rect -4384 6019 8664 6023
rect 8830 6132 18232 6137
rect 8830 6019 13856 6132
rect -4384 6014 13856 6019
rect 14022 6028 18232 6132
rect 18398 6057 23435 6146
rect 23601 6144 45246 6175
rect 23601 6057 27857 6144
rect 18398 6028 27857 6057
rect 14022 6026 27857 6028
rect 28023 6142 45246 6144
rect 28023 6141 35754 6142
rect 28023 6026 33030 6141
rect 14022 6023 33030 6026
rect 33196 6024 35754 6141
rect 35920 6024 45246 6142
rect 33196 6023 45246 6024
rect 14022 6014 45246 6023
rect -4384 5920 45246 6014
rect 46070 5920 46513 6288
rect -4384 5902 46513 5920
rect -5587 5881 46513 5902
rect -5587 5880 43159 5881
rect 44792 5880 46513 5881
rect -9849 5207 -1751 5224
rect 48849 5219 51439 7507
rect 42805 5207 51439 5219
rect -9849 4995 51439 5207
rect -9849 4900 2173 4995
rect 2310 4994 51439 4995
rect 2310 4991 31065 4994
rect 2310 4990 11745 4991
rect 2310 4900 6872 4990
rect -9849 4895 6872 4900
rect 7009 4896 11745 4990
rect 11882 4986 31065 4991
rect 11882 4985 26261 4986
rect 11882 4984 21381 4985
rect 11882 4896 16561 4984
rect 7009 4895 16561 4896
rect -9849 4889 16561 4895
rect 16698 4890 21381 4984
rect 21518 4891 26261 4985
rect 26398 4899 31065 4986
rect 31202 4990 51439 4994
rect 31202 4899 37116 4990
rect 26398 4895 37116 4899
rect 37253 4895 51439 4990
rect 26398 4891 51439 4895
rect 21518 4890 51439 4891
rect 16698 4889 51439 4890
rect -9849 4761 51439 4889
rect -9849 2363 -7261 4761
rect -3120 4760 51439 4761
rect -3120 4756 -2305 4760
rect 42805 4756 51439 4760
rect 42988 3529 46521 3531
rect 42808 3527 46521 3529
rect -2352 3525 46521 3527
rect -5738 3505 46521 3525
rect -5738 3098 -5349 3505
rect -4498 3499 46521 3505
rect -4498 3368 45192 3499
rect -4498 3358 35753 3368
rect -4498 3357 18226 3358
rect -4498 3352 8657 3357
rect -4498 3234 364 3352
rect 530 3339 8657 3352
rect 530 3234 3837 3339
rect -4498 3221 3837 3234
rect 4003 3239 8657 3339
rect 8823 3354 18226 3357
rect 8823 3239 13858 3354
rect 4003 3236 13858 3239
rect 14024 3240 18226 3354
rect 18392 3332 35753 3358
rect 18392 3330 33004 3332
rect 18392 3240 23433 3330
rect 14024 3236 23433 3240
rect 4003 3221 23433 3236
rect -4498 3212 23433 3221
rect 23599 3321 33004 3330
rect 23599 3212 27873 3321
rect -4498 3203 27873 3212
rect 28039 3214 33004 3321
rect 33170 3250 35753 3332
rect 35919 3250 45192 3368
rect 33170 3214 45192 3250
rect 28039 3203 45192 3214
rect -4498 3119 45192 3203
rect 46104 3119 46521 3499
rect -4498 3098 46521 3119
rect -5738 3080 46521 3098
rect 42808 3079 46521 3080
rect -9849 2351 -1481 2363
rect 48849 2362 51439 4756
rect 42835 2351 51439 2362
rect -9849 2197 51439 2351
rect -9849 2191 31069 2197
rect -9849 2190 11748 2191
rect -9849 2187 6874 2190
rect -9849 2092 2171 2187
rect 2308 2095 6874 2187
rect 7011 2096 11748 2190
rect 11885 2190 31069 2191
rect 11885 2096 16565 2190
rect 7011 2095 16565 2096
rect 16702 2188 31069 2190
rect 16702 2186 26252 2188
rect 16702 2095 21382 2186
rect 2308 2092 21382 2095
rect -9849 2091 21382 2092
rect 21519 2093 26252 2186
rect 26389 2102 31069 2188
rect 31206 2151 51439 2197
rect 31206 2102 37117 2151
rect 26389 2093 37117 2102
rect 21519 2091 37117 2093
rect -9849 2056 37117 2091
rect 37254 2056 51439 2151
rect -9849 1904 51439 2056
rect -9849 1900 -1481 1904
rect -9849 -212 -7261 1900
rect 42835 1899 51439 1904
rect -5687 671 -1817 677
rect 42691 671 46592 675
rect -5687 663 46592 671
rect -5687 653 45293 663
rect -5687 246 -5047 653
rect -4196 502 45293 653
rect -4196 489 3831 502
rect -4196 371 359 489
rect 525 384 3831 489
rect 3997 501 45293 502
rect 3997 499 23406 501
rect 3997 484 18221 499
rect 3997 483 13863 484
rect 3997 384 8648 483
rect 525 371 8648 384
rect -4196 365 8648 371
rect 8814 366 13863 483
rect 14029 381 18221 484
rect 18387 383 23406 499
rect 23572 492 45293 501
rect 23572 474 33018 492
rect 23572 383 27873 474
rect 18387 381 27873 383
rect 14029 366 27873 381
rect 8814 365 27873 366
rect -4196 356 27873 365
rect 28039 374 33018 474
rect 33184 374 35762 492
rect 35928 374 45293 492
rect 28039 356 45293 374
rect -4196 246 45293 356
rect -5687 245 45293 246
rect 46226 245 46592 663
rect -5687 225 46592 245
rect -5687 224 43159 225
rect -5687 219 -1817 224
rect 42863 223 43159 224
rect 48849 -212 51439 1899
rect -9849 -327 51439 -212
rect -9849 -393 16535 -327
rect -9849 -402 11709 -393
rect -9849 -657 2128 -402
rect 2367 -431 11709 -402
rect 2367 -657 6823 -431
rect -9849 -696 6823 -657
rect 7082 -606 11709 -431
rect 11938 -602 16535 -393
rect 16756 -368 51439 -327
rect 16756 -380 37051 -368
rect 16756 -414 26205 -380
rect 16756 -602 21332 -414
rect 11938 -606 21332 -602
rect 7082 -664 21332 -606
rect 21563 -637 26205 -414
rect 26428 -393 37051 -380
rect 26428 -637 31011 -393
rect 21563 -662 31011 -637
rect 31255 -659 37051 -393
rect 37326 -659 51439 -368
rect 31255 -662 51439 -659
rect 21563 -664 51439 -662
rect 7082 -696 51439 -664
rect -9849 -812 51439 -696
rect -9849 -5151 -7261 -812
rect 2069 -5151 2405 -812
rect 6761 -5151 7140 -812
rect 11630 -5151 12009 -812
rect 16442 -5151 16821 -812
rect 21293 -5151 21672 -812
rect 26111 -5151 26490 -812
rect -9852 -5152 26764 -5151
rect -9852 -5153 29998 -5152
rect 30968 -5153 31347 -812
rect 36993 -5153 37372 -812
rect 48849 -3734 51439 -812
rect 48851 -5153 51439 -3734
rect -9852 -7740 51444 -5153
rect -9852 -7745 -6438 -7740
rect 29811 -7741 51444 -7740
use 4MSB_weighted_binary  4MSB_weighted_binary_0
timestamp 1755845627
transform -1 0 43958 0 1 26320
box 2352 -4032 10080 56
use 6MSB_MATRIX  6MSB_MATRIX_0
timestamp 1755162181
transform 1 0 -2298 0 1 21392
box 2298 -21392 43904 2632
<< labels >>
flabel metal2 33432 26544 33768 26880 1 FreeSans 3200 0 0 0 X2
port 2 nsew signal input
flabel metal2 31920 26544 32256 26880 1 FreeSans 3200 0 0 0 X3
port 3 nsew signal input
flabel metal2 30184 26544 30520 26880 1 FreeSans 3200 0 0 0 X4
port 4 nsew signal input
flabel metal2 25536 26544 25872 26880 1 FreeSans 3200 0 0 0 X5
port 5 nsew signal input
flabel metal2 21840 26544 22176 26880 1 FreeSans 3200 0 0 0 X6
port 6 nsew signal input
flabel metal3 17192 26544 17528 26880 1 FreeSans 3200 0 0 0 X7
port 7 nsew signal input
flabel metal1 11424 26544 11760 26880 1 FreeSans 3200 0 0 0 X8
port 8 nsew signal input
flabel metal2 8344 26544 8680 26880 1 FreeSans 3200 0 0 0 X9
port 9 nsew signal input
flabel metal3 3415 26543 3752 26881 1 FreeSans 3200 0 0 0 X10
port 10 nsew signal input
flabel metal3 40264 26376 40600 26712 1 FreeSans 3200 0 0 0 VBIAS
port 13 nsew power bidirectional
flabel metal2 40768 27047 41104 27383 1 FreeSans 3200 0 0 0 OUTP
port 11 nsew power bidirectional
flabel metal2 35168 26880 35504 27216 1 FreeSans 3200 0 0 0 X1
port 1 nsew signal input
flabel metal2 38920 26320 39256 26656 1 FreeSans 3200 0 0 0 CLK
port 14 nsew signal bidirectional
rlabel metal4 27800 -3594 46988 -1006 1 VDD
port 15 n
rlabel metal4 -6204 -3592 -3615 30196 1 VDD
port 15 n
rlabel metal4 -6204 -3592 -312 -1009 1 VDD
port 15 n
flabel space -9852 32223 51436 34811 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel space 48851 -5153 51436 32223 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel space -9852 -7745 51444 -5153 1 FreeSans 8000 0 0 0 VSS
port 16 n
flabel space -9849 -5153 -7264 32223 1 FreeSans 8000 0 0 0 VSS
port 16 n
rlabel space 44397 -3597 46985 30190 1 VDD
port 15 n
rlabel metal4 -2581 -3591 27907 -1002 1 VDD
port 15 n
flabel metal4 -1571 27719 41443 30193 1 FreeSans 8000 0 0 0 VDD
port 15 nsew power bidirectional
rlabel metal4 -6209 27719 44816 30193 1 VDD
port 15 n
flabel metal3 3163 35114 3983 35941 1 FreeSans 6400 0 0 0 X10
port 10 n
flabel metal2 8112 35100 8932 35927 1 FreeSans 6400 0 0 0 X9
port 9 n
flabel metal2 11159 35023 11979 35850 1 FreeSans 6400 0 0 0 X8
port 8 n
flabel metal3 16944 35100 17764 35927 1 FreeSans 6400 0 0 0 X7
port 7 n
flabel metal2 21602 35265 22422 36092 1 FreeSans 6400 0 0 0 X6
port 6 n
flabel metal2 25299 35318 26119 36145 1 FreeSans 6400 0 0 0 X5
port 5 n
flabel metal2 29980 35246 30800 36073 1 FreeSans 6400 0 0 0 X4
port 4 n
flabel metal2 31704 35276 32524 36103 1 FreeSans 6400 0 0 0 X3
port 3 n
flabel metal2 33185 35283 34005 36110 1 FreeSans 6400 0 0 0 X2
port 2 n
flabel metal2 34937 35280 35757 36107 1 FreeSans 6400 0 0 0 X1
port 1 n
flabel metal2 38668 35091 39488 35918 1 FreeSans 6400 0 0 0 CLK
port 14 n
flabel metal2 41269 26040 41608 26376 1 FreeSans 3200 0 0 0 OUTN
port 12 nsew power bidirectional
flabel metal3 40053 36415 40873 37242 1 FreeSans 6400 1 0 0 VBIAS
port 13 n
flabel metal2 51734 26958 52331 27523 1 FreeSans 6400 1 0 0 OUTP
port 11 n
flabel metal2 52349 25424 52946 25989 1 FreeSans 6400 1 0 0 OUTN
port 12 n
<< end >>
