magic
tech gf180mcuD
magscale 1 10
timestamp 1755923713
<< nwell >>
rect 18259 -970 18308 -918
rect 3478 -6067 3590 -5601
rect 4037 -5666 4089 -5614
rect 2863 -11970 2929 -11959
rect 37953 -14068 38013 -14012
<< pwell >>
rect 3478 -5601 3590 -5163
<< mvpmos >>
rect 2863 -11970 2929 -11959
<< polysilicon >>
rect 37955 -2868 38011 -2815
rect 4037 -5666 4089 -5614
<< metal1 >>
rect 2800 2497 37912 2632
rect 2800 2494 28000 2497
rect 2800 2492 13496 2494
rect 2800 2436 3696 2492
rect 3752 2436 8568 2492
rect 8624 2438 13496 2492
rect 13552 2492 28000 2494
rect 13552 2491 23184 2492
rect 13552 2438 18256 2491
rect 8624 2436 18256 2438
rect 2800 2435 18256 2436
rect 18312 2436 23184 2491
rect 23240 2441 28000 2492
rect 28056 2464 37912 2497
rect 28056 2441 32872 2464
rect 23240 2436 32872 2441
rect 18312 2435 32872 2436
rect 2800 2408 32872 2435
rect 32928 2408 37744 2464
rect 37800 2408 37912 2464
rect 2800 2296 37912 2408
rect 11997 1323 12498 1400
rect 13020 1361 13787 1438
rect 3483 1195 6151 1315
rect 13710 1273 13787 1361
rect 17975 1343 18634 1421
rect 21615 1383 22231 1457
rect 22722 1387 23474 1461
rect 13710 1206 13719 1273
rect 13776 1206 13787 1273
rect 13710 1181 13787 1206
rect 18556 1254 18634 1343
rect 18556 1188 18565 1254
rect 18626 1188 18634 1254
rect 23399 1298 23474 1387
rect 27799 1334 28354 1417
rect 31308 1380 31922 1470
rect 32432 1350 33173 1440
rect 23399 1229 23407 1298
rect 23464 1229 23474 1298
rect 23399 1192 23474 1229
rect 28268 1287 28354 1334
rect 28268 1224 28280 1287
rect 28337 1224 28354 1287
rect 28268 1196 28354 1224
rect 33082 1262 33173 1350
rect 33082 1202 33095 1262
rect 33156 1202 33173 1262
rect 18556 1166 18634 1188
rect 33082 1179 33173 1202
rect 3099 805 4095 870
rect 4028 537 4095 805
rect 43568 672 43904 1400
rect 4028 485 4032 537
rect 4088 485 4095 537
rect 8008 504 43904 672
rect 4028 472 4095 485
rect 3487 291 3714 411
rect 4812 84 5370 103
rect 4437 80 5370 84
rect 4406 39 5370 80
rect 4406 37 4852 39
rect 4406 16 4437 37
rect 4929 -73 5485 -9
rect 3494 -613 3805 -373
rect 4929 -576 4993 -73
rect 3681 -983 3700 -907
rect 3768 -983 3807 -907
rect 8040 -965 8116 504
rect 9658 91 10300 103
rect 9283 82 10300 91
rect 9212 39 10300 82
rect 9212 37 9698 39
rect 9212 18 9283 37
rect 9775 -73 10705 -9
rect 8872 -280 8944 -127
rect 9775 -387 9839 -73
rect 8559 -983 8574 -907
rect 8632 -983 8738 -907
rect 12886 -965 12962 504
rect 14504 91 15146 103
rect 14058 39 15146 91
rect 14058 37 14544 39
rect 14058 27 14129 37
rect 14621 -73 15551 -9
rect 13718 -188 13790 -152
rect 14621 -613 14685 -73
rect 17732 -965 17808 504
rect 19350 90 19992 103
rect 18904 39 19992 90
rect 18904 37 19390 39
rect 18904 26 18975 37
rect 19467 -73 20397 -9
rect 19467 -613 19531 -73
rect 18247 -918 18359 -907
rect 18247 -970 18259 -918
rect 18311 -970 18359 -918
rect 22578 -965 22654 504
rect 24196 94 24838 103
rect 23750 39 24838 94
rect 23750 37 24236 39
rect 23750 30 23821 37
rect 24313 -73 25243 -9
rect 24313 -613 24377 -73
rect 27424 -965 27500 504
rect 29042 93 29684 103
rect 28596 39 29684 93
rect 28596 37 29082 39
rect 28596 29 28667 37
rect 29159 -73 30089 -9
rect 29159 -613 29223 -73
rect 27978 -918 28083 -907
rect 18247 -983 18359 -970
rect 27978 -971 28001 -918
rect 28056 -971 28083 -918
rect 32270 -965 32346 504
rect 33888 93 34530 103
rect 33442 39 34530 93
rect 33442 37 33928 39
rect 33442 29 33513 37
rect 34005 -73 34935 -9
rect 33102 -183 33174 -153
rect 34005 -613 34069 -73
rect 32849 -915 32941 -907
rect 27978 -983 28083 -971
rect 32849 -972 32869 -915
rect 32932 -972 32941 -915
rect 37116 -965 37192 504
rect 37746 148 37796 340
rect 38734 95 39376 103
rect 38287 39 39376 95
rect 38287 37 38773 39
rect 38287 31 38359 37
rect 38851 -73 39781 -9
rect 38851 -613 38915 -73
rect 41962 -965 42038 504
rect 32849 -983 32941 -972
rect 3511 -1397 3753 -1277
rect 43568 -2128 43904 504
rect 8008 -2296 43904 -2128
rect 4846 -2700 5484 -2697
rect 4846 -2756 4896 -2700
rect 4952 -2756 5484 -2700
rect 4846 -2761 5484 -2756
rect 4406 -2873 5280 -2809
rect 3499 -3413 3749 -3293
rect 3671 -3783 3687 -3707
rect 3755 -3783 3835 -3707
rect 8040 -3765 8116 -2296
rect 9713 -2701 10374 -2697
rect 9713 -2757 9775 -2701
rect 9831 -2757 10374 -2701
rect 9713 -2761 10374 -2757
rect 9230 -2873 10144 -2809
rect 8549 -3783 8568 -3707
rect 8628 -3783 8728 -3707
rect 12886 -3765 12962 -2296
rect 14549 -2701 15056 -2697
rect 14549 -2757 14584 -2701
rect 14640 -2757 15056 -2701
rect 14549 -2761 15056 -2757
rect 14093 -2873 15025 -2809
rect 17732 -3765 17808 -2296
rect 19371 -2701 19899 -2697
rect 19371 -2757 19460 -2701
rect 19516 -2757 19899 -2701
rect 19371 -2761 19899 -2757
rect 18905 -2873 20398 -2809
rect 18248 -3719 18368 -3707
rect 18248 -3773 18261 -3719
rect 18319 -3773 18368 -3719
rect 22578 -3765 22654 -2296
rect 24212 -2700 24784 -2697
rect 24212 -2756 24273 -2700
rect 24329 -2756 24784 -2700
rect 24212 -2761 24784 -2756
rect 23789 -2873 25283 -2809
rect 18248 -3783 18368 -3773
rect 27424 -3765 27500 -2296
rect 29050 -2699 29560 -2697
rect 29050 -2755 29147 -2699
rect 29203 -2755 29560 -2699
rect 29050 -2761 29560 -2755
rect 28617 -2873 30052 -2809
rect 27980 -3718 28079 -3707
rect 27980 -3770 27993 -3718
rect 28049 -3770 28079 -3718
rect 32270 -3765 32346 -2296
rect 33926 -2701 34786 -2697
rect 33926 -2757 33993 -2701
rect 34049 -2757 34786 -2701
rect 33926 -2761 34786 -2757
rect 33465 -2873 34789 -2809
rect 32854 -3714 32935 -3707
rect 27980 -3783 28079 -3770
rect 32854 -3774 32869 -3714
rect 32932 -3774 32935 -3714
rect 37116 -3765 37192 -2296
rect 37746 -2652 37796 -2492
rect 38769 -2699 39440 -2697
rect 38769 -2755 38835 -2699
rect 38891 -2755 39440 -2699
rect 38769 -2761 39440 -2755
rect 38350 -2873 39689 -2809
rect 41962 -3765 42038 -2296
rect 32854 -3783 32935 -3774
rect 3496 -4197 3720 -4077
rect 43568 -4928 43904 -2296
rect 8008 -5096 43904 -4928
rect 3370 -5309 3709 -5189
rect 4846 -5500 5484 -5497
rect 4846 -5556 4896 -5500
rect 4952 -5556 5484 -5500
rect 4846 -5561 5484 -5556
rect 4406 -5673 5280 -5609
rect 3294 -6213 3701 -5973
rect 3678 -6583 3691 -6507
rect 3750 -6583 3829 -6507
rect 8040 -6565 8116 -5096
rect 9713 -5499 10374 -5497
rect 9713 -5555 9775 -5499
rect 9831 -5555 10374 -5499
rect 9713 -5561 10374 -5555
rect 9230 -5673 10144 -5609
rect 8548 -6583 8565 -6507
rect 8624 -6583 8714 -6507
rect 12886 -6565 12962 -5096
rect 14549 -5501 15056 -5497
rect 14549 -5557 14584 -5501
rect 14640 -5557 15056 -5501
rect 14549 -5561 15056 -5557
rect 14093 -5673 15025 -5609
rect 17732 -6565 17808 -5096
rect 19371 -5501 19899 -5497
rect 19371 -5557 19461 -5501
rect 19517 -5557 19899 -5501
rect 19371 -5561 19899 -5557
rect 18905 -5673 20398 -5609
rect 18246 -6520 18369 -6507
rect 18246 -6573 18257 -6520
rect 18315 -6573 18369 -6520
rect 22578 -6565 22654 -5096
rect 24212 -5502 24784 -5497
rect 24212 -5558 24273 -5502
rect 24329 -5558 24784 -5502
rect 24212 -5561 24784 -5558
rect 23789 -5673 25283 -5609
rect 27424 -6565 27500 -5096
rect 29050 -5502 29560 -5497
rect 29050 -5558 29147 -5502
rect 29203 -5558 29560 -5502
rect 29050 -5561 29560 -5558
rect 28617 -5673 30052 -5609
rect 27973 -6519 28070 -6507
rect 18246 -6583 18369 -6573
rect 27973 -6574 27989 -6519
rect 28042 -6574 28070 -6519
rect 32270 -6565 32346 -5096
rect 33926 -5502 34767 -5497
rect 33926 -5558 33992 -5502
rect 34048 -5558 34767 -5502
rect 33926 -5561 34767 -5558
rect 33465 -5673 34789 -5609
rect 32858 -6518 32939 -6507
rect 27973 -6583 28070 -6574
rect 32858 -6573 32870 -6518
rect 32933 -6573 32939 -6518
rect 37116 -6565 37192 -5096
rect 37745 -5452 37796 -5284
rect 38769 -5506 39440 -5497
rect 38769 -5558 38833 -5506
rect 38894 -5558 39440 -5506
rect 38769 -5561 39440 -5558
rect 38350 -5673 39689 -5609
rect 41962 -6565 42038 -5096
rect 32858 -6583 32939 -6573
rect 3454 -6997 3459 -6877
rect 3468 -6997 3793 -6877
rect 42521 -7728 42924 -7727
rect 43568 -7728 43904 -5096
rect 8008 -7896 43904 -7728
rect 4846 -8301 5484 -8297
rect 4846 -8357 4895 -8301
rect 4951 -8357 5484 -8301
rect 4846 -8361 5484 -8357
rect 4406 -8473 5280 -8409
rect 3493 -9013 3697 -8893
rect 3656 -9317 3851 -9307
rect 3656 -9373 3696 -9317
rect 3752 -9373 3851 -9317
rect 8040 -9365 8116 -7896
rect 9713 -8302 10374 -8297
rect 9713 -8358 9775 -8302
rect 9831 -8358 10374 -8302
rect 9713 -8361 10374 -8358
rect 9230 -8473 10144 -8409
rect 3656 -9383 3851 -9373
rect 8551 -9383 8566 -9307
rect 8627 -9383 8704 -9307
rect 12886 -9365 12962 -7896
rect 14549 -8302 15056 -8297
rect 14549 -8358 14584 -8302
rect 14640 -8358 15056 -8302
rect 14549 -8361 15056 -8358
rect 14093 -8473 15025 -8409
rect 17732 -9365 17808 -7896
rect 19371 -8301 19899 -8297
rect 19371 -8357 19460 -8301
rect 19516 -8357 19899 -8301
rect 19371 -8361 19899 -8357
rect 18905 -8473 20398 -8409
rect 18241 -9321 18368 -9307
rect 18241 -9373 18256 -9321
rect 18314 -9373 18368 -9321
rect 22578 -9365 22654 -7896
rect 24212 -8301 24784 -8297
rect 24212 -8357 24273 -8301
rect 24329 -8357 24784 -8301
rect 24212 -8361 24784 -8357
rect 23789 -8473 25283 -8409
rect 27424 -9365 27500 -7896
rect 29050 -8302 29560 -8297
rect 29050 -8358 29148 -8302
rect 29204 -8358 29560 -8302
rect 29050 -8361 29560 -8358
rect 28617 -8473 30052 -8409
rect 27976 -9317 28074 -9307
rect 18241 -9383 18368 -9373
rect 27976 -9375 27993 -9317
rect 28053 -9375 28074 -9317
rect 32270 -9365 32346 -7896
rect 33926 -8302 34713 -8297
rect 33926 -8358 33992 -8302
rect 34048 -8358 34713 -8302
rect 33926 -8361 34713 -8358
rect 33465 -8473 34789 -8409
rect 32853 -9317 32953 -9307
rect 27976 -9383 28074 -9375
rect 32853 -9372 32868 -9317
rect 32932 -9372 32953 -9317
rect 37116 -9365 37192 -7896
rect 37745 -8252 37796 -8092
rect 38769 -8301 39440 -8297
rect 38769 -8357 38835 -8301
rect 38891 -8357 39440 -8301
rect 38769 -8361 39440 -8357
rect 38350 -8473 39689 -8409
rect 41962 -9365 42038 -7896
rect 32853 -9383 32953 -9372
rect 3491 -9797 3708 -9677
rect 43568 -10528 43904 -7896
rect 8008 -10696 43904 -10528
rect 3489 -10909 3772 -10789
rect 4846 -11100 5484 -11097
rect 4846 -11156 4895 -11100
rect 4951 -11156 5484 -11100
rect 4846 -11161 5484 -11156
rect 4406 -11273 5280 -11209
rect 3513 -11574 3818 -11573
rect 3505 -11693 3818 -11574
rect 3499 -11813 3818 -11693
rect 2863 -11970 2929 -11959
rect 3676 -12183 3688 -12107
rect 3758 -12183 3872 -12107
rect 8040 -12165 8116 -10696
rect 9713 -11101 10374 -11097
rect 9713 -11157 9776 -11101
rect 9832 -11157 10374 -11101
rect 9713 -11161 10374 -11157
rect 9230 -11273 10144 -11209
rect 8541 -12118 8702 -12107
rect 8541 -12171 8562 -12118
rect 8614 -12171 8702 -12118
rect 12886 -12165 12962 -10696
rect 14549 -11102 15056 -11097
rect 14549 -11158 14586 -11102
rect 14642 -11158 15056 -11102
rect 14549 -11161 15056 -11158
rect 14093 -11273 15025 -11209
rect 17732 -12165 17808 -10696
rect 19371 -11099 19899 -11097
rect 19371 -11155 19461 -11099
rect 19517 -11155 19899 -11099
rect 19371 -11161 19899 -11155
rect 18905 -11273 20398 -11209
rect 18239 -12121 18373 -12107
rect 8541 -12183 8702 -12171
rect 18239 -12174 18253 -12121
rect 18309 -12174 18373 -12121
rect 22578 -12165 22654 -10696
rect 24212 -11100 24784 -11097
rect 24212 -11156 24274 -11100
rect 24330 -11156 24784 -11100
rect 24212 -11161 24784 -11156
rect 23789 -11273 25283 -11209
rect 27424 -12165 27500 -10696
rect 29050 -11100 29560 -11097
rect 29050 -11156 29148 -11100
rect 29204 -11156 29560 -11100
rect 29050 -11161 29560 -11156
rect 28617 -11273 30052 -11209
rect 27983 -12117 28075 -12107
rect 18239 -12183 18373 -12174
rect 27983 -12175 27998 -12117
rect 28058 -12175 28075 -12117
rect 32270 -12165 32346 -10696
rect 33926 -11099 34788 -11097
rect 33926 -11155 33993 -11099
rect 34049 -11155 34788 -11099
rect 33926 -11161 34788 -11155
rect 33465 -11273 34789 -11209
rect 32836 -12119 32933 -12107
rect 27983 -12183 28075 -12175
rect 32836 -12171 32889 -12119
rect 37116 -12165 37192 -10696
rect 37744 -11052 37796 -10893
rect 38769 -11100 39440 -11097
rect 38769 -11156 38835 -11100
rect 38891 -11156 39440 -11100
rect 38769 -11161 39440 -11156
rect 38350 -11273 39689 -11209
rect 41962 -12165 42038 -10696
rect 32836 -12183 32933 -12171
rect 3501 -12597 3765 -12477
rect 42537 -13328 42916 -13327
rect 43568 -13328 43904 -10696
rect 8008 -13496 9762 -13328
rect 9844 -13496 14570 -13328
rect 14655 -13496 24259 -13328
rect 24344 -13496 43904 -13328
rect 4846 -13902 5484 -13897
rect 4846 -13958 4895 -13902
rect 4951 -13958 5484 -13902
rect 4846 -13961 5484 -13958
rect 4406 -14073 5280 -14009
rect 3498 -14613 3710 -14493
rect 3668 -14983 3681 -14907
rect 3746 -14983 3864 -14907
rect 8040 -14965 8116 -13496
rect 9713 -13901 10374 -13897
rect 9713 -13957 9775 -13901
rect 9831 -13957 10374 -13901
rect 9713 -13961 10374 -13957
rect 9230 -14073 10144 -14009
rect 8561 -14919 8697 -14907
rect 8561 -14971 8581 -14919
rect 8633 -14971 8697 -14919
rect 12886 -14965 12962 -13496
rect 14549 -13902 15056 -13897
rect 14549 -13958 14585 -13902
rect 14641 -13958 15056 -13902
rect 14549 -13961 15056 -13958
rect 14093 -14073 15025 -14009
rect 17732 -14965 17808 -13496
rect 19371 -13900 19899 -13897
rect 19371 -13956 19462 -13900
rect 19518 -13956 19899 -13900
rect 19371 -13961 19899 -13956
rect 18905 -14073 20398 -14009
rect 18243 -14921 18383 -14907
rect 8561 -14983 8697 -14971
rect 18243 -14974 18256 -14921
rect 18312 -14974 18383 -14921
rect 22578 -14965 22654 -13496
rect 24212 -13901 24784 -13897
rect 24212 -13957 24274 -13901
rect 24330 -13957 24784 -13901
rect 24212 -13961 24784 -13957
rect 23789 -14073 25283 -14009
rect 27424 -14965 27500 -13496
rect 29050 -13900 29560 -13897
rect 29050 -13956 29147 -13900
rect 29203 -13956 29560 -13900
rect 29050 -13961 29560 -13956
rect 28617 -14073 30052 -14009
rect 27977 -14916 28064 -14907
rect 18243 -14983 18383 -14974
rect 27977 -14972 27997 -14916
rect 28062 -14972 28064 -14916
rect 32270 -14965 32346 -13496
rect 33926 -13900 34722 -13897
rect 33926 -13956 33991 -13900
rect 34047 -13956 34722 -13900
rect 33926 -13961 34722 -13956
rect 33465 -14073 34789 -14009
rect 32847 -14918 32968 -14907
rect 27977 -14983 28064 -14972
rect 32847 -14973 32868 -14918
rect 32936 -14973 32968 -14918
rect 37116 -14965 37192 -13496
rect 37751 -13709 37796 -13704
rect 37750 -13852 37796 -13709
rect 38769 -13901 39440 -13897
rect 38769 -13957 38835 -13901
rect 38891 -13957 39440 -13901
rect 38769 -13961 39440 -13957
rect 38350 -14073 39689 -14009
rect 41962 -14965 42038 -13496
rect 32847 -14983 32968 -14973
rect 3485 -15397 3712 -15277
rect 43568 -16128 43904 -13496
rect 8008 -16296 43904 -16128
rect 3473 -16509 3739 -16389
rect 4846 -16700 5484 -16697
rect 4846 -16756 4897 -16700
rect 4953 -16756 5484 -16700
rect 4846 -16761 5484 -16756
rect 4406 -16873 5280 -16809
rect 3455 -17413 3462 -17173
rect 3486 -17413 3722 -17173
rect 3674 -17783 3692 -17707
rect 3760 -17783 3881 -17707
rect 8040 -17765 8116 -16296
rect 9713 -16700 10374 -16697
rect 9713 -16756 9775 -16700
rect 9831 -16756 10374 -16700
rect 9713 -16761 10374 -16756
rect 9230 -16873 10144 -16809
rect 8551 -17720 8709 -17707
rect 8551 -17772 8572 -17720
rect 8626 -17772 8709 -17720
rect 12886 -17765 12962 -16296
rect 14549 -16701 15056 -16697
rect 14549 -16757 14585 -16701
rect 14641 -16757 15056 -16701
rect 14549 -16761 15056 -16757
rect 14093 -16873 15025 -16809
rect 17732 -17765 17808 -16296
rect 19371 -16701 19899 -16697
rect 19371 -16757 19462 -16701
rect 19518 -16757 19899 -16701
rect 19371 -16761 19899 -16757
rect 18905 -16873 20398 -16809
rect 18239 -17717 18381 -17707
rect 8551 -17783 8709 -17772
rect 18239 -17773 18253 -17717
rect 18315 -17773 18381 -17717
rect 22578 -17765 22654 -16296
rect 24212 -16702 24784 -16697
rect 24212 -16758 24274 -16702
rect 24330 -16758 24784 -16702
rect 24212 -16761 24784 -16758
rect 23789 -16873 25283 -16809
rect 18239 -17783 18381 -17773
rect 27424 -17765 27500 -16296
rect 29050 -16702 29560 -16697
rect 29050 -16758 29148 -16702
rect 29204 -16758 29560 -16702
rect 29050 -16761 29560 -16758
rect 28617 -16873 30052 -16809
rect 27987 -17716 28062 -17707
rect 27987 -17769 27999 -17716
rect 28060 -17769 28062 -17716
rect 32270 -17765 32346 -16296
rect 33926 -16700 34695 -16697
rect 33926 -16756 33993 -16700
rect 34049 -16756 34695 -16700
rect 33926 -16761 34695 -16756
rect 33465 -16873 34789 -16809
rect 32842 -17715 32947 -17707
rect 27987 -17783 28062 -17769
rect 32842 -17775 32868 -17715
rect 32935 -17775 32947 -17715
rect 37116 -17765 37192 -16296
rect 37748 -16652 37796 -16486
rect 38769 -16701 39440 -16697
rect 38769 -16757 38835 -16701
rect 38891 -16757 39440 -16701
rect 38769 -16761 39440 -16757
rect 38350 -16873 39689 -16809
rect 41962 -17765 42038 -16296
rect 32842 -17783 32947 -17775
rect 3492 -18197 3695 -18077
rect 38732 -18928 38984 -18927
rect 43568 -18928 43904 -16296
rect 8008 -19096 43904 -18928
rect 3824 -19452 3874 -19286
rect 4846 -19502 5484 -19497
rect 4846 -19555 4893 -19502
rect 4956 -19555 5484 -19502
rect 4846 -19561 5484 -19555
rect 4406 -19673 5280 -19609
rect 3679 -20583 3696 -20507
rect 3752 -20583 3853 -20507
rect 8040 -20565 8116 -19096
rect 8670 -19452 8720 -19286
rect 9713 -19501 10374 -19497
rect 9713 -19554 9772 -19501
rect 9834 -19554 10374 -19501
rect 9713 -19561 10374 -19554
rect 9230 -19673 10144 -19609
rect 8557 -20518 8706 -20507
rect 8557 -20570 8568 -20518
rect 8620 -20570 8706 -20518
rect 12886 -20565 12962 -19096
rect 13516 -19452 13566 -19286
rect 14549 -19505 15056 -19497
rect 14549 -19557 14580 -19505
rect 14645 -19557 15056 -19505
rect 14549 -19561 15056 -19557
rect 14093 -19673 15025 -19609
rect 17732 -20565 17808 -19096
rect 18362 -19452 18412 -19286
rect 19371 -19506 19899 -19497
rect 19371 -19558 19458 -19506
rect 19521 -19558 19899 -19506
rect 19371 -19561 19899 -19558
rect 18905 -19673 20398 -19609
rect 18239 -20521 18374 -20507
rect 8557 -20583 8706 -20570
rect 18239 -20577 18254 -20521
rect 18312 -20577 18374 -20521
rect 22578 -20565 22654 -19096
rect 23208 -19452 23258 -19286
rect 24212 -19503 24784 -19497
rect 24212 -19556 24269 -19503
rect 24334 -19556 24784 -19503
rect 24212 -19561 24784 -19556
rect 23789 -19673 25283 -19609
rect 27424 -20565 27500 -19096
rect 28054 -19452 28104 -19286
rect 29050 -19505 29560 -19497
rect 29050 -19558 29145 -19505
rect 29206 -19558 29560 -19505
rect 29050 -19561 29560 -19558
rect 28617 -19673 30052 -19609
rect 27988 -20517 28074 -20507
rect 27988 -20574 27998 -20517
rect 28059 -20574 28074 -20517
rect 32270 -20565 32346 -19096
rect 32900 -19452 32950 -19286
rect 33926 -19505 35419 -19497
rect 33926 -19557 33989 -19505
rect 34051 -19557 35419 -19505
rect 33926 -19561 35419 -19557
rect 33465 -19673 34789 -19609
rect 32844 -20517 32953 -20507
rect 18239 -20583 18374 -20577
rect 27988 -20583 28074 -20574
rect 32844 -20574 32869 -20517
rect 32932 -20574 32953 -20517
rect 37116 -20565 37192 -19096
rect 43568 -19219 43904 -19096
rect 32844 -20583 32953 -20574
<< via1 >>
rect 3696 2436 3752 2492
rect 8568 2436 8624 2492
rect 13496 2438 13552 2494
rect 18256 2435 18312 2491
rect 23184 2436 23240 2492
rect 28000 2441 28056 2497
rect 32872 2408 32928 2464
rect 37744 2408 37800 2464
rect 3107 1757 3167 1818
rect 13719 1206 13776 1273
rect 18565 1188 18626 1254
rect 23407 1229 23464 1298
rect 28280 1224 28337 1287
rect 33095 1202 33156 1262
rect 2765 836 2823 890
rect 6722 822 6785 883
rect 4032 485 4088 537
rect 3811 -11 3871 48
rect 4035 -67 4089 -15
rect 3107 -314 3167 -197
rect 2769 -776 2822 -683
rect 3099 -993 3170 -937
rect 3700 -983 3768 -907
rect 7569 -952 7623 -899
rect 8648 -88 8720 -36
rect 8882 -66 8934 -14
rect 8574 -983 8632 -907
rect 12415 -952 12469 -899
rect 13502 -90 13558 -34
rect 13727 -67 13782 -15
rect 13505 -974 13567 -916
rect 17261 -952 17315 -899
rect 18340 -91 18412 -39
rect 18573 -68 18628 -15
rect 18259 -970 18311 -918
rect 22107 -952 22161 -899
rect 23194 -10 23249 42
rect 23420 -67 23474 -14
rect 23199 -968 23256 -916
rect 26953 -952 27007 -899
rect 28040 -11 28094 42
rect 28264 -67 28322 -15
rect 28001 -971 28056 -918
rect 31799 -952 31853 -899
rect 32887 -9 32940 43
rect 33111 -68 33166 -15
rect 32869 -972 32932 -915
rect 36645 -952 36699 -899
rect 37957 -67 38013 -12
rect 37744 -971 37800 -915
rect 41491 -952 41545 -899
rect 7602 -1104 7656 -1051
rect 8019 -1103 8073 -1050
rect 12448 -1104 12502 -1051
rect 12865 -1103 12919 -1050
rect 17294 -1104 17348 -1051
rect 17711 -1103 17765 -1050
rect 22140 -1104 22194 -1051
rect 22557 -1103 22611 -1050
rect 26986 -1104 27040 -1051
rect 27403 -1103 27457 -1050
rect 31832 -1104 31886 -1051
rect 32249 -1103 32303 -1050
rect 36678 -1104 36732 -1051
rect 37095 -1103 37149 -1050
rect 41524 -1104 41578 -1051
rect 41941 -1103 41995 -1050
rect 4896 -2756 4952 -2700
rect 3812 -2811 3866 -2757
rect 4037 -2867 4090 -2814
rect 3092 -3790 3148 -3734
rect 3687 -3783 3755 -3707
rect 7569 -3752 7623 -3699
rect 8657 -2811 8712 -2756
rect 9775 -2757 9831 -2701
rect 8882 -2867 8936 -2815
rect 8568 -3783 8628 -3707
rect 12415 -3752 12469 -3699
rect 14584 -2757 14640 -2701
rect 13503 -2810 13559 -2758
rect 13727 -2867 13782 -2814
rect 13510 -3772 13566 -3717
rect 17261 -3752 17315 -3699
rect 18348 -2811 18403 -2754
rect 19460 -2757 19516 -2701
rect 18573 -2867 18627 -2815
rect 18261 -3773 18319 -3719
rect 22107 -3752 22161 -3699
rect 24273 -2756 24329 -2700
rect 23195 -2810 23249 -2758
rect 23418 -2868 23472 -2815
rect 23194 -3774 23253 -3718
rect 26953 -3752 27007 -3699
rect 29147 -2755 29203 -2699
rect 28041 -2810 28094 -2758
rect 28267 -2866 28320 -2812
rect 27993 -3770 28049 -3718
rect 31799 -3752 31853 -3699
rect 33993 -2757 34049 -2701
rect 32887 -2811 32941 -2757
rect 33112 -2867 33164 -2815
rect 32869 -3774 32932 -3714
rect 36645 -3752 36699 -3699
rect 38835 -2755 38891 -2699
rect 37955 -2868 38011 -2815
rect 37744 -3770 37800 -3714
rect 41491 -3752 41545 -3699
rect 7602 -3904 7656 -3851
rect 8019 -3903 8073 -3850
rect 12448 -3904 12502 -3851
rect 12865 -3903 12919 -3850
rect 17294 -3904 17348 -3851
rect 17711 -3903 17765 -3850
rect 22140 -3904 22194 -3851
rect 22557 -3903 22611 -3850
rect 26986 -3904 27040 -3851
rect 27403 -3903 27457 -3850
rect 31832 -3904 31886 -3851
rect 32249 -3903 32303 -3850
rect 36678 -3904 36732 -3851
rect 37095 -3903 37149 -3850
rect 41524 -3904 41578 -3851
rect 41941 -3903 41995 -3850
rect 3811 -5611 3867 -5555
rect 4896 -5556 4952 -5500
rect 4037 -5666 4089 -5614
rect 3076 -5907 3146 -5826
rect 2750 -6351 2803 -6277
rect 3087 -6592 3143 -6536
rect 3691 -6583 3750 -6507
rect 7569 -6552 7623 -6499
rect 9775 -5555 9831 -5499
rect 8656 -5611 8712 -5555
rect 8882 -5667 8935 -5615
rect 8565 -6583 8624 -6507
rect 12415 -6552 12469 -6499
rect 14584 -5557 14640 -5501
rect 13500 -5611 13563 -5558
rect 13728 -5667 13780 -5615
rect 13508 -6571 13566 -6515
rect 17261 -6552 17315 -6499
rect 19461 -5557 19517 -5501
rect 18350 -5610 18409 -5557
rect 18574 -5667 18629 -5612
rect 18257 -6573 18315 -6520
rect 22107 -6552 22161 -6499
rect 23190 -5608 23251 -5556
rect 24273 -5558 24329 -5502
rect 23420 -5667 23473 -5614
rect 23194 -6572 23250 -6517
rect 26953 -6552 27007 -6499
rect 29147 -5558 29203 -5502
rect 28041 -5611 28098 -5559
rect 28267 -5666 28319 -5614
rect 27989 -6574 28042 -6519
rect 31799 -6552 31853 -6499
rect 33992 -5558 34048 -5502
rect 32887 -5611 32945 -5559
rect 33111 -5667 33165 -5614
rect 32870 -6573 32933 -6518
rect 36645 -6552 36699 -6499
rect 38833 -5558 38894 -5506
rect 37956 -5667 38012 -5612
rect 37744 -6570 37800 -6514
rect 41491 -6552 41545 -6499
rect 7602 -6704 7656 -6651
rect 8019 -6703 8073 -6650
rect 12448 -6704 12502 -6651
rect 12865 -6703 12919 -6650
rect 17294 -6704 17348 -6651
rect 17711 -6703 17765 -6650
rect 22140 -6704 22194 -6651
rect 22557 -6703 22611 -6650
rect 26986 -6704 27040 -6651
rect 27403 -6703 27457 -6650
rect 31832 -6704 31886 -6651
rect 32249 -6703 32303 -6650
rect 36678 -6704 36732 -6651
rect 37095 -6703 37149 -6650
rect 41524 -6704 41578 -6651
rect 41941 -6703 41995 -6650
rect 3810 -8412 3868 -8356
rect 4895 -8357 4951 -8301
rect 4036 -8467 4089 -8415
rect 3696 -9373 3752 -9317
rect 7569 -9352 7623 -9299
rect 9775 -8358 9831 -8302
rect 8656 -8411 8714 -8358
rect 8882 -8469 8938 -8414
rect 8566 -9383 8627 -9307
rect 12415 -9352 12469 -9299
rect 14584 -8358 14640 -8302
rect 13500 -8411 13561 -8359
rect 13728 -8467 13780 -8415
rect 13510 -9371 13567 -9316
rect 17261 -9352 17315 -9299
rect 19460 -8357 19516 -8301
rect 18347 -8412 18407 -8357
rect 18571 -8470 18629 -8412
rect 18256 -9373 18314 -9321
rect 22107 -9352 22161 -9299
rect 24273 -8357 24329 -8301
rect 23196 -8411 23251 -8359
rect 23420 -8468 23475 -8413
rect 23196 -9371 23250 -9316
rect 26953 -9352 27007 -9299
rect 28042 -8409 28097 -8357
rect 29148 -8358 29204 -8302
rect 28264 -8467 28321 -8413
rect 27993 -9375 28053 -9317
rect 31799 -9352 31853 -9299
rect 33992 -8358 34048 -8302
rect 32886 -8413 32943 -8360
rect 33110 -8469 33165 -8414
rect 32868 -9372 32932 -9317
rect 36645 -9352 36699 -9299
rect 38835 -8357 38891 -8301
rect 37957 -8467 38012 -8414
rect 37744 -9371 37800 -9315
rect 41491 -9352 41545 -9299
rect 3302 -9439 3358 -9383
rect 7602 -9504 7656 -9451
rect 8019 -9503 8073 -9450
rect 12448 -9504 12502 -9451
rect 12865 -9503 12919 -9450
rect 17294 -9504 17348 -9451
rect 17711 -9503 17765 -9450
rect 22140 -9504 22194 -9451
rect 22557 -9503 22611 -9450
rect 26986 -9504 27040 -9451
rect 27403 -9503 27457 -9450
rect 31832 -9504 31886 -9451
rect 32249 -9503 32303 -9450
rect 36678 -9504 36732 -9451
rect 37095 -9503 37149 -9450
rect 41524 -9504 41578 -9451
rect 41941 -9503 41995 -9450
rect 4895 -11156 4951 -11100
rect 3811 -11292 3867 -11236
rect 4037 -11266 4089 -11214
rect 3096 -11514 3157 -11421
rect 2865 -11959 2926 -11876
rect 3203 -12225 3259 -12169
rect 3688 -12183 3758 -12107
rect 7569 -12152 7623 -12099
rect 8654 -11212 8710 -11156
rect 9776 -11157 9832 -11101
rect 8874 -11272 8938 -11212
rect 8562 -12171 8614 -12118
rect 12415 -12152 12469 -12099
rect 14586 -11158 14642 -11102
rect 13502 -11210 13557 -11158
rect 13728 -11266 13780 -11214
rect 13506 -12171 13560 -12119
rect 17261 -12152 17315 -12099
rect 19461 -11155 19517 -11099
rect 18347 -11209 18404 -11155
rect 18573 -11268 18626 -11213
rect 18253 -12174 18309 -12121
rect 22107 -12152 22161 -12099
rect 24274 -11156 24330 -11100
rect 23194 -11208 23253 -11156
rect 23420 -11267 23477 -11213
rect 23192 -12173 23252 -12116
rect 26953 -12152 27007 -12099
rect 29148 -11156 29204 -11100
rect 28039 -11212 28098 -11158
rect 28266 -11266 28318 -11214
rect 27998 -12175 28058 -12117
rect 31799 -12152 31853 -12099
rect 33993 -11155 34049 -11099
rect 32888 -11211 32947 -11156
rect 33111 -11268 33164 -11216
rect 32889 -12171 32941 -12119
rect 36645 -12152 36699 -12099
rect 38835 -11156 38891 -11100
rect 37957 -11268 38013 -11212
rect 37744 -12170 37800 -12114
rect 41491 -12152 41545 -12099
rect 7602 -12304 7656 -12251
rect 8019 -12303 8073 -12250
rect 12448 -12304 12502 -12251
rect 12865 -12303 12919 -12250
rect 17294 -12304 17348 -12251
rect 17711 -12303 17765 -12250
rect 22140 -12304 22194 -12251
rect 22557 -12303 22611 -12250
rect 26986 -12304 27040 -12251
rect 27403 -12303 27457 -12250
rect 31832 -12304 31886 -12251
rect 32249 -12303 32303 -12250
rect 36678 -12304 36732 -12251
rect 37095 -12303 37149 -12250
rect 41524 -12304 41578 -12251
rect 41941 -12303 41995 -12250
rect 4895 -13958 4951 -13902
rect 3808 -14088 3871 -14035
rect 4037 -14067 4089 -14015
rect 3187 -14963 3243 -14907
rect 3681 -14983 3746 -14907
rect 7569 -14952 7623 -14899
rect 9775 -13957 9831 -13901
rect 8657 -14012 8712 -13957
rect 8882 -14067 8937 -14013
rect 8581 -14971 8633 -14919
rect 12415 -14952 12469 -14899
rect 13504 -14010 13559 -13956
rect 14585 -13958 14641 -13902
rect 13727 -14067 13782 -14014
rect 13512 -14971 13567 -14918
rect 17261 -14952 17315 -14899
rect 18348 -14011 18406 -13955
rect 19462 -13956 19518 -13900
rect 18572 -14068 18630 -14013
rect 18256 -14974 18312 -14921
rect 22107 -14952 22161 -14899
rect 24274 -13957 24330 -13901
rect 23196 -14011 23255 -13957
rect 23419 -14068 23474 -14015
rect 23196 -14971 23251 -14913
rect 26953 -14952 27007 -14899
rect 28039 -14012 28099 -13950
rect 29147 -13956 29203 -13900
rect 28264 -14067 28320 -14013
rect 27997 -14972 28062 -14916
rect 31799 -14952 31853 -14899
rect 32885 -14014 32947 -13955
rect 33991 -13956 34047 -13900
rect 33112 -14067 33164 -14014
rect 32868 -14973 32936 -14918
rect 36645 -14952 36699 -14899
rect 38835 -13957 38891 -13901
rect 37957 -14067 38013 -14013
rect 37744 -14970 37800 -14914
rect 41491 -14952 41545 -14899
rect 7602 -15104 7656 -15051
rect 8019 -15103 8073 -15050
rect 12448 -15104 12502 -15051
rect 12865 -15103 12919 -15050
rect 17294 -15104 17348 -15051
rect 17711 -15103 17765 -15050
rect 22140 -15104 22194 -15051
rect 22557 -15103 22611 -15050
rect 26986 -15104 27040 -15051
rect 27403 -15103 27457 -15050
rect 31832 -15104 31886 -15051
rect 32249 -15103 32303 -15050
rect 36678 -15104 36732 -15051
rect 37095 -15103 37149 -15050
rect 41524 -15104 41578 -15051
rect 41941 -15103 41995 -15050
rect 4897 -16756 4953 -16700
rect 3181 -16883 3251 -16806
rect 3809 -16891 3865 -16835
rect 4036 -16867 4088 -16815
rect 2850 -17778 2911 -17716
rect 3692 -17783 3760 -17707
rect 7569 -17752 7623 -17699
rect 9775 -16756 9831 -16700
rect 8654 -16811 8713 -16757
rect 8882 -16867 8934 -16815
rect 8572 -17772 8626 -17720
rect 12415 -17752 12469 -17699
rect 13501 -16811 13560 -16754
rect 14585 -16757 14641 -16701
rect 13728 -16867 13783 -16814
rect 13507 -17769 13559 -17717
rect 17261 -17752 17315 -17699
rect 19462 -16757 19518 -16701
rect 18346 -16815 18407 -16758
rect 18573 -16868 18627 -16814
rect 18253 -17773 18315 -17717
rect 22107 -17752 22161 -17699
rect 23194 -16811 23252 -16757
rect 24274 -16758 24330 -16702
rect 23419 -16867 23475 -16814
rect 23197 -17775 23250 -17714
rect 26953 -17752 27007 -17699
rect 28037 -16811 28101 -16754
rect 29148 -16758 29204 -16702
rect 28267 -16866 28320 -16814
rect 27999 -17769 28060 -17716
rect 31799 -17752 31853 -17699
rect 32884 -16811 32943 -16755
rect 33993 -16756 34049 -16700
rect 33112 -16867 33165 -16815
rect 32868 -17775 32935 -17715
rect 36645 -17752 36699 -17699
rect 38835 -16757 38891 -16701
rect 37952 -16870 38016 -16812
rect 37744 -17772 37800 -17716
rect 41491 -17752 41545 -17699
rect 7602 -17904 7656 -17851
rect 8019 -17903 8073 -17850
rect 12448 -17904 12502 -17851
rect 12865 -17903 12919 -17850
rect 17294 -17904 17348 -17851
rect 17711 -17903 17765 -17850
rect 22140 -17904 22194 -17851
rect 22557 -17903 22611 -17850
rect 26986 -17904 27040 -17851
rect 27403 -17903 27457 -17850
rect 31832 -17904 31886 -17851
rect 32249 -17903 32303 -17850
rect 36678 -17904 36732 -17851
rect 37095 -17903 37149 -17850
rect 41524 -17904 41578 -17851
rect 41941 -17903 41995 -17850
rect 4893 -19555 4956 -19502
rect 4036 -19668 4089 -19615
rect 3696 -20583 3752 -20507
rect 7569 -20552 7623 -20499
rect 9772 -19554 9834 -19501
rect 8882 -19666 8936 -19614
rect 8568 -20570 8620 -20518
rect 12415 -20552 12469 -20499
rect 14580 -19557 14645 -19505
rect 13729 -19666 13781 -19614
rect 13515 -20570 13568 -20518
rect 17261 -20552 17315 -20499
rect 19458 -19558 19521 -19506
rect 18573 -19669 18630 -19613
rect 18254 -20577 18312 -20521
rect 22107 -20552 22161 -20499
rect 24269 -19556 24334 -19503
rect 23419 -19667 23474 -19615
rect 23198 -20574 23250 -20517
rect 26953 -20552 27007 -20499
rect 29145 -19558 29206 -19505
rect 28263 -19667 28318 -19614
rect 27998 -20574 28059 -20517
rect 31799 -20552 31853 -20499
rect 33989 -19557 34051 -19505
rect 33111 -19668 33166 -19614
rect 32869 -20574 32932 -20517
rect 36645 -20552 36699 -20499
rect 7602 -20704 7656 -20651
rect 8019 -20703 8073 -20650
rect 12448 -20704 12502 -20651
rect 12865 -20703 12919 -20650
rect 17294 -20704 17348 -20651
rect 17711 -20703 17765 -20650
rect 22140 -20704 22194 -20651
rect 22557 -20703 22611 -20650
rect 26986 -20704 27040 -20651
rect 27403 -20703 27457 -20650
rect 31832 -20704 31886 -20651
rect 32249 -20703 32303 -20650
rect 36678 -20704 36732 -20651
rect 37095 -20703 37149 -20650
<< metal2 >>
rect 3686 2492 3762 2502
rect 3686 2436 3696 2492
rect 3752 2436 3762 2492
rect 3686 2426 3762 2436
rect 8558 2492 8634 2502
rect 8558 2436 8568 2492
rect 8624 2436 8634 2492
rect 8558 2426 8634 2436
rect 13486 2494 13562 2504
rect 13486 2438 13496 2494
rect 13552 2438 13562 2494
rect 13486 2428 13562 2438
rect 18246 2491 18322 2501
rect 18246 2435 18256 2491
rect 18312 2435 18322 2491
rect 18246 2425 18322 2435
rect 23174 2492 23250 2502
rect 23174 2436 23184 2492
rect 23240 2436 23250 2492
rect 23174 2426 23250 2436
rect 27987 2497 28069 2509
rect 27987 2441 28000 2497
rect 28056 2441 28069 2497
rect 27987 2429 28069 2441
rect 32858 2464 32939 2476
rect 32858 2408 32872 2464
rect 32928 2408 32939 2464
rect 32858 2394 32939 2408
rect 37734 2464 37810 2474
rect 37734 2408 37744 2464
rect 37800 2408 37810 2464
rect 37734 2398 37810 2408
rect 3089 1818 3185 1835
rect 3089 1757 3107 1818
rect 3167 1757 3185 1818
rect 3089 1736 3185 1757
rect 2749 890 2835 897
rect 2749 836 2765 890
rect 2823 889 2835 890
rect 3101 889 3169 1736
rect 23370 1301 23497 1314
rect 13688 1278 13804 1299
rect 13688 1203 13716 1278
rect 13780 1203 13804 1278
rect 13688 1181 13804 1203
rect 18536 1257 18648 1264
rect 18536 1185 18562 1257
rect 18631 1185 18648 1257
rect 23370 1223 23403 1301
rect 23468 1223 23497 1301
rect 23370 1196 23497 1223
rect 28247 1291 28370 1304
rect 28247 1218 28271 1291
rect 28344 1218 28370 1291
rect 28247 1192 28370 1218
rect 33065 1262 33188 1274
rect 33065 1202 33095 1262
rect 33156 1202 33188 1262
rect 18536 1166 18648 1185
rect 33065 1176 33188 1202
rect 43064 896 43400 1400
rect 2823 836 3170 889
rect 2749 821 3170 836
rect 6693 888 6807 894
rect 6693 819 6718 888
rect 6790 819 6807 888
rect 6693 804 6807 819
rect 7504 728 43400 896
rect 3998 537 4115 539
rect 3998 480 4029 537
rect 4093 480 4115 537
rect 3998 448 4115 480
rect 3798 53 3887 57
rect 3509 48 3887 53
rect 3509 -11 3811 48
rect 3871 -11 3887 48
rect 3509 -13 3887 -11
rect 3099 -197 3170 -163
rect 3099 -255 3107 -197
rect 2759 -314 3107 -255
rect 3167 -314 3170 -197
rect 2759 -327 3170 -314
rect 2759 -683 2831 -327
rect 2759 -776 2769 -683
rect 2822 -776 2831 -683
rect 2759 -800 2831 -776
rect 3089 -937 3183 -928
rect 3089 -993 3099 -937
rect 3170 -993 3183 -937
rect 3089 -1002 3183 -993
rect 3099 -1736 3170 -1002
rect 3099 -1820 3170 -1792
rect 3509 -1722 3585 -13
rect 3798 -22 3887 -13
rect 4010 -13 4115 -1
rect 4010 -69 4033 -13
rect 4092 -69 4115 -13
rect 4010 -78 4115 -69
rect 3672 -907 3794 -884
rect 3672 -983 3696 -907
rect 3774 -983 3794 -907
rect 7558 -899 7634 728
rect 8859 -12 8951 -8
rect 7558 -952 7569 -899
rect 7623 -952 7634 -899
rect 7558 -965 7634 -952
rect 8391 -36 8768 -27
rect 8391 -88 8648 -36
rect 8720 -88 8768 -36
rect 8859 -68 8880 -12
rect 8938 -68 8951 -12
rect 8859 -74 8951 -68
rect 8391 -103 8768 -88
rect 3672 -1002 3794 -983
rect 7591 -1050 8083 -1039
rect 7591 -1051 8019 -1050
rect 7591 -1104 7602 -1051
rect 7656 -1103 8019 -1051
rect 8073 -1103 8083 -1050
rect 7656 -1104 8083 -1103
rect 7591 -1115 8083 -1104
rect 7798 -1456 7874 -1115
rect 8391 -1334 8467 -103
rect 8545 -907 8658 -893
rect 8545 -983 8574 -907
rect 8632 -983 8658 -907
rect 12404 -899 12480 728
rect 13701 -13 13810 -1
rect 12404 -952 12415 -899
rect 12469 -952 12480 -899
rect 12404 -965 12480 -952
rect 13262 -34 13608 -31
rect 13262 -90 13502 -34
rect 13558 -90 13608 -34
rect 13701 -69 13725 -13
rect 13784 -69 13810 -13
rect 13701 -78 13810 -69
rect 13262 -104 13608 -90
rect 8545 -1000 8658 -983
rect 12437 -1050 12929 -1039
rect 12437 -1051 12865 -1050
rect 12437 -1104 12448 -1051
rect 12502 -1103 12865 -1051
rect 12919 -1103 12929 -1050
rect 12502 -1104 12929 -1103
rect 12437 -1115 12929 -1104
rect 8391 -1400 8467 -1390
rect 12644 -1456 12720 -1115
rect 13262 -1333 13338 -104
rect 13469 -916 13581 -896
rect 13469 -974 13505 -916
rect 13567 -974 13581 -916
rect 17250 -899 17326 728
rect 18553 -12 18646 2
rect 17250 -952 17261 -899
rect 17315 -952 17326 -899
rect 17250 -965 17326 -952
rect 18079 -39 18464 -29
rect 18079 -91 18340 -39
rect 18412 -91 18464 -39
rect 18553 -70 18570 -12
rect 18632 -70 18646 -12
rect 18553 -84 18646 -70
rect 18079 -105 18464 -91
rect 13469 -998 13581 -974
rect 17283 -1050 17775 -1039
rect 17283 -1051 17711 -1050
rect 17283 -1104 17294 -1051
rect 17348 -1103 17711 -1051
rect 17765 -1103 17775 -1050
rect 17348 -1104 17775 -1103
rect 17283 -1115 17775 -1104
rect 13262 -1400 13338 -1389
rect 17490 -1456 17566 -1115
rect 18079 -1324 18157 -105
rect 18223 -915 18325 -896
rect 18223 -972 18256 -915
rect 18315 -972 18325 -915
rect 22096 -899 22172 728
rect 22953 42 23263 48
rect 22953 20 23194 42
rect 22096 -952 22107 -899
rect 22161 -952 22172 -899
rect 22096 -965 22172 -952
rect 22952 -10 23194 20
rect 23249 -10 23263 42
rect 22952 -16 23263 -10
rect 23405 -12 23487 -1
rect 18223 -996 18325 -972
rect 22129 -1050 22621 -1039
rect 22129 -1051 22557 -1050
rect 22129 -1104 22140 -1051
rect 22194 -1103 22557 -1051
rect 22611 -1103 22621 -1050
rect 22194 -1104 22621 -1103
rect 22129 -1115 22621 -1104
rect 18079 -1398 18157 -1380
rect 22336 -1456 22412 -1115
rect 22952 -1335 23028 -16
rect 23405 -69 23418 -12
rect 23476 -69 23487 -12
rect 23405 -80 23487 -69
rect 23156 -913 23270 -895
rect 23156 -971 23194 -913
rect 23260 -971 23270 -913
rect 26942 -899 27018 728
rect 26942 -952 26953 -899
rect 27007 -952 27018 -899
rect 26942 -965 27018 -952
rect 27766 42 28133 49
rect 27766 -11 28040 42
rect 28094 -11 28133 42
rect 27766 -22 28133 -11
rect 28249 -13 28338 1
rect 23156 -999 23270 -971
rect 26975 -1050 27467 -1039
rect 26975 -1051 27403 -1050
rect 26975 -1104 26986 -1051
rect 27040 -1103 27403 -1051
rect 27457 -1103 27467 -1050
rect 27040 -1104 27467 -1103
rect 26975 -1115 27467 -1104
rect 22952 -1391 22962 -1335
rect 23018 -1391 23028 -1335
rect 22952 -1400 23028 -1391
rect 27182 -1456 27258 -1115
rect 27766 -1334 27842 -22
rect 28249 -69 28262 -13
rect 28325 -69 28338 -13
rect 28249 -83 28338 -69
rect 27975 -915 28081 -898
rect 27975 -975 27999 -915
rect 28058 -975 28081 -915
rect 31788 -899 31864 728
rect 31788 -952 31799 -899
rect 31853 -952 31864 -899
rect 31788 -965 31864 -952
rect 32637 43 32964 47
rect 32637 -9 32887 43
rect 32940 -9 32964 43
rect 32637 -13 32964 -9
rect 33097 -13 33182 -3
rect 27975 -1001 28081 -975
rect 31821 -1050 32313 -1039
rect 31821 -1051 32249 -1050
rect 31821 -1104 31832 -1051
rect 31886 -1103 32249 -1051
rect 32303 -1103 32313 -1050
rect 31886 -1104 32313 -1103
rect 31821 -1115 32313 -1104
rect 27766 -1390 27778 -1334
rect 27834 -1390 27842 -1334
rect 27766 -1400 27842 -1390
rect 32028 -1456 32104 -1115
rect 32637 -1336 32713 -13
rect 33097 -70 33109 -13
rect 33168 -70 33182 -13
rect 33097 -79 33182 -70
rect 32850 -915 32947 -897
rect 32850 -972 32869 -915
rect 32932 -972 32947 -915
rect 36634 -899 36710 728
rect 36634 -952 36645 -899
rect 36699 -952 36710 -899
rect 36634 -965 36710 -952
rect 37482 -12 38026 -3
rect 37482 -67 37957 -12
rect 38013 -67 38026 -12
rect 37482 -80 38026 -67
rect 32850 -990 32947 -972
rect 36667 -1050 37159 -1039
rect 36667 -1051 37095 -1050
rect 36667 -1104 36678 -1051
rect 36732 -1103 37095 -1051
rect 37149 -1103 37159 -1050
rect 36732 -1104 37159 -1103
rect 36667 -1115 37159 -1104
rect 32637 -1392 32647 -1336
rect 32703 -1392 32713 -1336
rect 32637 -1400 32713 -1392
rect 36874 -1456 36950 -1115
rect 37482 -1335 37558 -80
rect 41480 -899 41556 728
rect 37732 -915 37811 -905
rect 37732 -971 37744 -915
rect 37800 -971 37811 -915
rect 41480 -952 41491 -899
rect 41545 -952 41556 -899
rect 41480 -965 41556 -952
rect 37732 -981 37811 -971
rect 41513 -1050 42005 -1039
rect 41513 -1051 41941 -1050
rect 41513 -1104 41524 -1051
rect 41578 -1103 41941 -1051
rect 41995 -1103 42005 -1050
rect 41578 -1104 42005 -1103
rect 41513 -1115 42005 -1104
rect 37482 -1391 37492 -1335
rect 37548 -1391 37558 -1335
rect 37482 -1400 37558 -1391
rect 41720 -1456 41796 -1115
rect 7392 -1512 42881 -1456
rect 7392 -1568 42672 -1512
rect 42728 -1568 42881 -1512
rect 7392 -1624 42881 -1568
rect 3509 -1788 3514 -1722
rect 3582 -1788 3585 -1722
rect 3509 -1818 3585 -1788
rect 4883 -1742 4966 -1680
rect 4883 -1798 4895 -1742
rect 4951 -1798 4966 -1742
rect 4883 -2700 4966 -1798
rect 43064 -1904 43400 728
rect 7504 -2072 43400 -1904
rect 3462 -2757 3903 -2745
rect 3462 -2811 3812 -2757
rect 3866 -2811 3903 -2757
rect 4883 -2756 4896 -2700
rect 4952 -2756 4966 -2700
rect 4883 -2761 4966 -2756
rect 3462 -2822 3903 -2811
rect 4009 -2812 4115 -2806
rect 3082 -3734 3158 -3707
rect 3082 -3790 3092 -3734
rect 3148 -3790 3158 -3734
rect 3082 -4551 3158 -3790
rect 3082 -4607 3092 -4551
rect 3148 -4607 3158 -4551
rect 3082 -4648 3158 -4607
rect 3462 -4538 3538 -2822
rect 4009 -2868 4035 -2812
rect 4092 -2868 4115 -2812
rect 4009 -2875 4115 -2868
rect 3655 -3707 3779 -3692
rect 3655 -3783 3687 -3707
rect 3755 -3783 3779 -3707
rect 7558 -3699 7634 -2072
rect 9762 -2136 9844 -2128
rect 9762 -2192 9776 -2136
rect 9832 -2192 9844 -2136
rect 9762 -2701 9844 -2192
rect 7558 -3752 7569 -3699
rect 7623 -3752 7634 -3699
rect 7558 -3765 7634 -3752
rect 8391 -2756 8742 -2749
rect 8391 -2811 8657 -2756
rect 8712 -2811 8742 -2756
rect 9762 -2757 9775 -2701
rect 9831 -2757 9844 -2701
rect 9762 -2761 9844 -2757
rect 8391 -2824 8742 -2811
rect 8860 -2812 8959 -2807
rect 3655 -3800 3779 -3783
rect 7591 -3850 8083 -3839
rect 7591 -3851 8019 -3850
rect 7591 -3904 7602 -3851
rect 7656 -3903 8019 -3851
rect 8073 -3903 8083 -3850
rect 7656 -3904 8083 -3903
rect 7591 -3915 8083 -3904
rect 7798 -4256 7874 -3915
rect 8391 -4131 8467 -2824
rect 8860 -2870 8879 -2812
rect 8938 -2870 8959 -2812
rect 8860 -2876 8959 -2870
rect 8539 -3707 8643 -3693
rect 8539 -3783 8568 -3707
rect 8628 -3783 8643 -3707
rect 12404 -3699 12480 -2072
rect 14570 -2137 14655 -2128
rect 14570 -2193 14584 -2137
rect 14640 -2193 14655 -2137
rect 14570 -2701 14655 -2193
rect 12404 -3752 12415 -3699
rect 12469 -3752 12480 -3699
rect 12404 -3765 12480 -3752
rect 13261 -2758 13595 -2749
rect 13261 -2810 13503 -2758
rect 13559 -2810 13595 -2758
rect 14570 -2757 14584 -2701
rect 14640 -2757 14655 -2701
rect 14570 -2760 14655 -2757
rect 13261 -2826 13595 -2810
rect 13704 -2812 13805 -2804
rect 8539 -3797 8643 -3783
rect 12437 -3850 12929 -3839
rect 12437 -3851 12865 -3850
rect 12437 -3904 12448 -3851
rect 12502 -3903 12865 -3851
rect 12919 -3903 12929 -3850
rect 12502 -3904 12929 -3903
rect 12437 -3915 12929 -3904
rect 8391 -4187 8401 -4131
rect 8457 -4187 8467 -4131
rect 8391 -4198 8467 -4187
rect 12644 -4256 12720 -3915
rect 13261 -4132 13337 -2826
rect 13704 -2869 13725 -2812
rect 13784 -2869 13805 -2812
rect 13704 -2882 13805 -2869
rect 13472 -3714 13586 -3692
rect 13472 -3774 13507 -3714
rect 13570 -3774 13586 -3714
rect 17250 -3699 17326 -2072
rect 19448 -2142 19531 -2134
rect 19448 -2198 19463 -2142
rect 19519 -2198 19531 -2142
rect 19448 -2701 19531 -2198
rect 17250 -3752 17261 -3699
rect 17315 -3752 17326 -3699
rect 17250 -3765 17326 -3752
rect 18080 -2754 18443 -2745
rect 18080 -2811 18348 -2754
rect 18403 -2811 18443 -2754
rect 19448 -2757 19460 -2701
rect 19516 -2757 19531 -2701
rect 19448 -2761 19531 -2757
rect 18080 -2823 18443 -2811
rect 18558 -2812 18642 -2798
rect 13472 -3803 13586 -3774
rect 17283 -3850 17775 -3839
rect 17283 -3851 17711 -3850
rect 17283 -3904 17294 -3851
rect 17348 -3903 17711 -3851
rect 17765 -3903 17775 -3850
rect 17348 -3904 17775 -3903
rect 17283 -3915 17775 -3904
rect 13261 -4188 13271 -4132
rect 13327 -4188 13337 -4132
rect 13261 -4200 13337 -4188
rect 17490 -4256 17566 -3915
rect 18080 -4122 18156 -2823
rect 18558 -2870 18570 -2812
rect 18629 -2870 18642 -2812
rect 18558 -2878 18642 -2870
rect 18233 -3716 18335 -3695
rect 18233 -3777 18259 -3716
rect 18323 -3777 18335 -3716
rect 22096 -3699 22172 -2072
rect 24259 -2139 24344 -2129
rect 24259 -2195 24273 -2139
rect 24329 -2195 24344 -2139
rect 24259 -2700 24344 -2195
rect 22096 -3752 22107 -3699
rect 22161 -3752 22172 -3699
rect 22096 -3765 22172 -3752
rect 22951 -2758 23271 -2754
rect 22951 -2810 23195 -2758
rect 23249 -2810 23271 -2758
rect 24259 -2756 24273 -2700
rect 24329 -2756 24344 -2700
rect 24259 -2761 24344 -2756
rect 22951 -2816 23271 -2810
rect 23402 -2813 23491 -2796
rect 18233 -3801 18335 -3777
rect 22129 -3850 22621 -3839
rect 22129 -3851 22557 -3850
rect 22129 -3904 22140 -3851
rect 22194 -3903 22557 -3851
rect 22611 -3903 22621 -3850
rect 22194 -3904 22621 -3903
rect 22129 -3915 22621 -3904
rect 18080 -4178 18090 -4122
rect 18146 -4178 18156 -4122
rect 18080 -4188 18156 -4178
rect 22336 -4256 22412 -3915
rect 22951 -4136 23027 -2816
rect 23402 -2870 23416 -2813
rect 23475 -2870 23491 -2813
rect 23402 -2883 23491 -2870
rect 26942 -3699 27018 -2072
rect 29135 -2140 29216 -2131
rect 29135 -2196 29147 -2140
rect 29203 -2196 29216 -2140
rect 29135 -2699 29216 -2196
rect 23155 -3718 23270 -3699
rect 23155 -3774 23194 -3718
rect 23253 -3774 23270 -3718
rect 26942 -3752 26953 -3699
rect 27007 -3752 27018 -3699
rect 26942 -3765 27018 -3752
rect 27767 -2758 28109 -2750
rect 27767 -2810 28041 -2758
rect 28094 -2810 28109 -2758
rect 29135 -2755 29147 -2699
rect 29203 -2755 29216 -2699
rect 29135 -2760 29216 -2755
rect 27767 -2817 28109 -2810
rect 28246 -2810 28340 -2801
rect 27767 -2905 27842 -2817
rect 28246 -2868 28265 -2810
rect 28322 -2868 28340 -2810
rect 28246 -2881 28340 -2868
rect 23155 -3796 23270 -3774
rect 26975 -3850 27467 -3839
rect 26975 -3851 27403 -3850
rect 26975 -3904 26986 -3851
rect 27040 -3903 27403 -3851
rect 27457 -3903 27467 -3850
rect 27040 -3904 27467 -3903
rect 26975 -3915 27467 -3904
rect 22951 -4192 22961 -4136
rect 23017 -4192 23027 -4136
rect 22951 -4200 23027 -4192
rect 27182 -4256 27258 -3915
rect 27767 -4135 27843 -2905
rect 27965 -3714 28068 -3696
rect 27965 -3772 27990 -3714
rect 28052 -3772 28068 -3714
rect 31788 -3699 31864 -2072
rect 33979 -2139 34061 -2129
rect 33979 -2195 33993 -2139
rect 34049 -2195 34061 -2139
rect 33979 -2701 34061 -2195
rect 31788 -3752 31799 -3699
rect 31853 -3752 31864 -3699
rect 31788 -3765 31864 -3752
rect 32639 -2757 32967 -2751
rect 32639 -2811 32887 -2757
rect 32941 -2811 32967 -2757
rect 33979 -2757 33993 -2701
rect 34049 -2757 34061 -2701
rect 33979 -2760 34061 -2757
rect 32639 -2819 32967 -2811
rect 33092 -2813 33180 -2801
rect 27965 -3796 28068 -3772
rect 31821 -3850 32313 -3839
rect 31821 -3851 32249 -3850
rect 31821 -3904 31832 -3851
rect 31886 -3903 32249 -3851
rect 32303 -3903 32313 -3850
rect 31886 -3904 32313 -3903
rect 31821 -3915 32313 -3904
rect 27767 -4191 27777 -4135
rect 27833 -4191 27843 -4135
rect 27767 -4200 27843 -4191
rect 32028 -4256 32104 -3915
rect 32639 -4135 32715 -2819
rect 33092 -2869 33110 -2813
rect 33166 -2869 33180 -2813
rect 33092 -2880 33180 -2869
rect 32843 -3714 32940 -3695
rect 32843 -3774 32869 -3714
rect 32932 -3774 32940 -3714
rect 36634 -3699 36710 -2072
rect 38823 -2139 38903 -2129
rect 38823 -2195 38835 -2139
rect 38891 -2195 38903 -2139
rect 38823 -2699 38903 -2195
rect 38823 -2755 38835 -2699
rect 38891 -2755 38903 -2699
rect 38823 -2757 38903 -2755
rect 36634 -3752 36645 -3699
rect 36699 -3752 36710 -3699
rect 36634 -3765 36710 -3752
rect 37455 -2815 38035 -2806
rect 37455 -2868 37955 -2815
rect 38011 -2868 38035 -2815
rect 37455 -2874 38035 -2868
rect 32843 -3788 32940 -3774
rect 36667 -3850 37159 -3839
rect 36667 -3851 37095 -3850
rect 36667 -3904 36678 -3851
rect 36732 -3903 37095 -3851
rect 37149 -3903 37159 -3850
rect 36732 -3904 37159 -3903
rect 36667 -3915 37159 -3904
rect 32639 -4191 32649 -4135
rect 32705 -4191 32715 -4135
rect 32639 -4200 32715 -4191
rect 36874 -4256 36950 -3915
rect 37455 -4136 37531 -2874
rect 41480 -3699 41556 -2072
rect 37731 -3714 37810 -3704
rect 37731 -3770 37744 -3714
rect 37800 -3770 37810 -3714
rect 41480 -3752 41491 -3699
rect 41545 -3752 41556 -3699
rect 41480 -3765 41556 -3752
rect 37731 -3780 37810 -3770
rect 41513 -3850 42005 -3839
rect 41513 -3851 41941 -3850
rect 41513 -3904 41524 -3851
rect 41578 -3903 41941 -3851
rect 41995 -3903 42005 -3850
rect 41578 -3904 42005 -3903
rect 41513 -3915 42005 -3904
rect 37455 -4192 37465 -4136
rect 37521 -4192 37531 -4136
rect 37455 -4200 37531 -4192
rect 41720 -4256 41796 -3915
rect 7392 -4312 42881 -4256
rect 7392 -4368 42672 -4312
rect 42728 -4368 42881 -4312
rect 7392 -4424 42881 -4368
rect 3462 -4594 3472 -4538
rect 3528 -4594 3538 -4538
rect 3462 -4648 3538 -4594
rect 4883 -4539 4966 -4480
rect 4883 -4595 4894 -4539
rect 4950 -4595 4966 -4539
rect 4883 -5500 4966 -4595
rect 43064 -4704 43400 -2072
rect 7504 -4872 43400 -4704
rect 3459 -5555 3890 -5544
rect 3459 -5611 3811 -5555
rect 3867 -5611 3890 -5555
rect 4883 -5556 4896 -5500
rect 4952 -5556 4966 -5500
rect 4883 -5560 4966 -5556
rect 3459 -5624 3890 -5611
rect 4015 -5612 4108 -5609
rect 3068 -5826 3150 -5773
rect 3068 -5840 3076 -5826
rect 2734 -5907 3076 -5840
rect 3146 -5907 3150 -5826
rect 2734 -5925 3150 -5907
rect 2734 -6277 2819 -5925
rect 2734 -6330 2750 -6277
rect 2740 -6351 2750 -6330
rect 2803 -6330 2819 -6277
rect 2803 -6351 2812 -6330
rect 2740 -6370 2812 -6351
rect 3077 -6536 3154 -6465
rect 3077 -6592 3087 -6536
rect 3143 -6592 3154 -6536
rect 3077 -7337 3154 -6592
rect 3077 -7393 3089 -7337
rect 3145 -7393 3154 -7337
rect 3077 -7448 3154 -7393
rect 3459 -7337 3535 -5624
rect 4015 -5668 4035 -5612
rect 4091 -5668 4108 -5612
rect 4015 -5675 4108 -5668
rect 3660 -6507 3762 -6493
rect 3660 -6583 3691 -6507
rect 3750 -6583 3762 -6507
rect 7558 -6499 7634 -4872
rect 9762 -4938 9844 -4928
rect 9762 -4994 9775 -4938
rect 9831 -4994 9844 -4938
rect 9762 -5499 9844 -4994
rect 7558 -6552 7569 -6499
rect 7623 -6552 7634 -6499
rect 7558 -6565 7634 -6552
rect 8389 -5555 8724 -5550
rect 8389 -5611 8656 -5555
rect 8712 -5611 8724 -5555
rect 9762 -5555 9775 -5499
rect 9831 -5555 9844 -5499
rect 9762 -5561 9844 -5555
rect 8389 -5622 8724 -5611
rect 8860 -5613 8955 -5608
rect 3660 -6600 3762 -6583
rect 7591 -6650 8083 -6639
rect 7591 -6651 8019 -6650
rect 7591 -6704 7602 -6651
rect 7656 -6703 8019 -6651
rect 8073 -6703 8083 -6650
rect 7656 -6704 8083 -6703
rect 7591 -6715 8083 -6704
rect 7798 -7056 7874 -6715
rect 8389 -6934 8465 -5622
rect 8860 -5670 8878 -5613
rect 8937 -5670 8955 -5613
rect 8860 -5674 8955 -5670
rect 8529 -6507 8634 -6496
rect 8529 -6583 8565 -6507
rect 8624 -6583 8634 -6507
rect 12404 -6499 12480 -4872
rect 14570 -4941 14655 -4928
rect 14570 -4997 14584 -4941
rect 14640 -4997 14655 -4941
rect 14570 -5501 14655 -4997
rect 12404 -6552 12415 -6499
rect 12469 -6552 12480 -6499
rect 12404 -6565 12480 -6552
rect 13240 -5558 13581 -5550
rect 13240 -5611 13500 -5558
rect 13563 -5611 13581 -5558
rect 14570 -5557 14584 -5501
rect 14640 -5557 14655 -5501
rect 14570 -5562 14655 -5557
rect 13240 -5619 13581 -5611
rect 13701 -5613 13802 -5602
rect 8529 -6597 8634 -6583
rect 12437 -6650 12929 -6639
rect 12437 -6651 12865 -6650
rect 12437 -6704 12448 -6651
rect 12502 -6703 12865 -6651
rect 12919 -6703 12929 -6650
rect 12502 -6704 12929 -6703
rect 12437 -6715 12929 -6704
rect 8389 -6990 8399 -6934
rect 8455 -6990 8465 -6934
rect 8389 -7000 8465 -6990
rect 12644 -7056 12720 -6715
rect 13240 -6926 13316 -5619
rect 13701 -5669 13725 -5613
rect 13783 -5669 13802 -5613
rect 13701 -5679 13802 -5669
rect 13470 -6513 13579 -6495
rect 13470 -6573 13506 -6513
rect 13569 -6573 13579 -6513
rect 17250 -6499 17326 -4872
rect 19448 -4937 19531 -4928
rect 19448 -4993 19462 -4937
rect 19518 -4993 19531 -4937
rect 19448 -5501 19531 -4993
rect 17250 -6552 17261 -6499
rect 17315 -6552 17326 -6499
rect 17250 -6565 17326 -6552
rect 18079 -5557 18425 -5553
rect 18079 -5610 18350 -5557
rect 18409 -5610 18425 -5557
rect 19448 -5557 19461 -5501
rect 19517 -5557 19531 -5501
rect 19448 -5562 19531 -5557
rect 18079 -5615 18425 -5610
rect 18556 -5607 18645 -5598
rect 13470 -6597 13579 -6573
rect 17283 -6650 17775 -6639
rect 17283 -6651 17711 -6650
rect 17283 -6704 17294 -6651
rect 17348 -6703 17711 -6651
rect 17765 -6703 17775 -6650
rect 17348 -6704 17775 -6703
rect 17283 -6715 17775 -6704
rect 13240 -6982 13250 -6926
rect 13306 -6982 13316 -6926
rect 13240 -6998 13316 -6982
rect 17490 -7056 17566 -6715
rect 18079 -6936 18155 -5615
rect 18556 -5671 18569 -5607
rect 18634 -5671 18645 -5607
rect 18556 -5682 18645 -5671
rect 18230 -6517 18333 -6492
rect 18230 -6577 18253 -6517
rect 18318 -6577 18333 -6517
rect 22096 -6499 22172 -4872
rect 24259 -4934 24344 -4928
rect 24259 -4990 24273 -4934
rect 24329 -4990 24344 -4934
rect 24259 -5502 24344 -4990
rect 22096 -6552 22107 -6499
rect 22161 -6552 22172 -6499
rect 22096 -6565 22172 -6552
rect 22950 -5556 23268 -5550
rect 22950 -5608 23190 -5556
rect 23251 -5608 23268 -5556
rect 24259 -5558 24273 -5502
rect 24329 -5558 24344 -5502
rect 24259 -5561 24344 -5558
rect 22950 -5616 23268 -5608
rect 23404 -5610 23490 -5601
rect 18230 -6599 18333 -6577
rect 22129 -6650 22621 -6639
rect 22129 -6651 22557 -6650
rect 22129 -6704 22140 -6651
rect 22194 -6703 22557 -6651
rect 22611 -6703 22621 -6650
rect 22194 -6704 22621 -6703
rect 22129 -6715 22621 -6704
rect 18079 -6992 18089 -6936
rect 18145 -6992 18155 -6936
rect 18079 -7000 18155 -6992
rect 22336 -7056 22412 -6715
rect 22950 -6937 23026 -5616
rect 23404 -5671 23416 -5610
rect 23478 -5671 23490 -5610
rect 23404 -5683 23490 -5671
rect 23153 -6516 23268 -6495
rect 23153 -6572 23194 -6516
rect 23252 -6572 23268 -6516
rect 26942 -6499 27018 -4872
rect 29135 -4935 29216 -4928
rect 29135 -4991 29147 -4935
rect 29203 -4991 29216 -4935
rect 29135 -5502 29216 -4991
rect 26942 -6552 26953 -6499
rect 27007 -6552 27018 -6499
rect 26942 -6565 27018 -6552
rect 27763 -5559 28113 -5545
rect 27763 -5611 28041 -5559
rect 28098 -5611 28113 -5559
rect 29135 -5558 29147 -5502
rect 29203 -5558 29216 -5502
rect 29135 -5561 29216 -5558
rect 27763 -5622 28113 -5611
rect 28251 -5611 28335 -5601
rect 23153 -6597 23268 -6572
rect 26975 -6650 27467 -6639
rect 26975 -6651 27403 -6650
rect 26975 -6704 26986 -6651
rect 27040 -6703 27403 -6651
rect 27457 -6703 27467 -6650
rect 27040 -6704 27467 -6703
rect 26975 -6715 27467 -6704
rect 22950 -6993 22960 -6937
rect 23016 -6993 23026 -6937
rect 22950 -7000 23026 -6993
rect 27182 -7056 27258 -6715
rect 27763 -6932 27839 -5622
rect 28251 -5668 28264 -5611
rect 28323 -5668 28335 -5611
rect 28251 -5683 28335 -5668
rect 27963 -6515 28073 -6494
rect 27963 -6576 27985 -6515
rect 28045 -6576 28073 -6515
rect 31788 -6499 31864 -4872
rect 33979 -4934 34061 -4928
rect 33979 -4990 33992 -4934
rect 34048 -4990 34061 -4934
rect 33979 -5502 34061 -4990
rect 31788 -6552 31799 -6499
rect 31853 -6552 31864 -6499
rect 31788 -6565 31864 -6552
rect 32639 -5559 32962 -5548
rect 32639 -5611 32887 -5559
rect 32945 -5611 32962 -5559
rect 33979 -5558 33992 -5502
rect 34048 -5558 34061 -5502
rect 33979 -5561 34061 -5558
rect 32639 -5626 32962 -5611
rect 33096 -5611 33179 -5606
rect 27963 -6597 28073 -6576
rect 31821 -6650 32313 -6639
rect 31821 -6651 32249 -6650
rect 31821 -6704 31832 -6651
rect 31886 -6703 32249 -6651
rect 32303 -6703 32313 -6650
rect 31886 -6704 32313 -6703
rect 31821 -6715 32313 -6704
rect 27763 -6988 27773 -6932
rect 27829 -6988 27839 -6932
rect 27763 -6996 27839 -6988
rect 32028 -7056 32104 -6715
rect 32639 -6934 32715 -5626
rect 33096 -5669 33109 -5611
rect 33169 -5669 33179 -5611
rect 33096 -5679 33179 -5669
rect 36634 -6499 36710 -4872
rect 38808 -5502 38920 -5497
rect 38808 -5558 38833 -5502
rect 38894 -5558 38920 -5502
rect 38808 -5561 38920 -5558
rect 32851 -6517 32944 -6500
rect 32851 -6573 32870 -6517
rect 32933 -6573 32944 -6517
rect 36634 -6552 36645 -6499
rect 36699 -6552 36710 -6499
rect 36634 -6565 36710 -6552
rect 37454 -5612 38029 -5602
rect 37454 -5667 37956 -5612
rect 38012 -5667 38029 -5612
rect 37454 -5679 38029 -5667
rect 32851 -6588 32944 -6573
rect 36667 -6650 37159 -6639
rect 36667 -6651 37095 -6650
rect 36667 -6704 36678 -6651
rect 36732 -6703 37095 -6651
rect 37149 -6703 37159 -6650
rect 36732 -6704 37159 -6703
rect 36667 -6715 37159 -6704
rect 32639 -6990 32649 -6934
rect 32705 -6990 32715 -6934
rect 32639 -6999 32715 -6990
rect 36874 -7056 36950 -6715
rect 37454 -7000 37530 -5679
rect 41480 -6499 41556 -4872
rect 37733 -6514 37811 -6503
rect 37733 -6570 37744 -6514
rect 37800 -6570 37811 -6514
rect 41480 -6552 41491 -6499
rect 41545 -6552 41556 -6499
rect 41480 -6565 41556 -6552
rect 37733 -6580 37811 -6570
rect 41513 -6650 42005 -6639
rect 41513 -6651 41941 -6650
rect 41513 -6704 41524 -6651
rect 41578 -6703 41941 -6651
rect 41995 -6703 42005 -6650
rect 41578 -6704 42005 -6703
rect 41513 -6715 42005 -6704
rect 41720 -7056 41796 -6715
rect 7392 -7112 42889 -7056
rect 7392 -7168 42671 -7112
rect 42728 -7168 42889 -7112
rect 7392 -7224 42889 -7168
rect 3459 -7393 3470 -7337
rect 3526 -7393 3535 -7337
rect 3459 -7448 3535 -7393
rect 4883 -7342 4966 -7280
rect 4883 -7398 4898 -7342
rect 4954 -7398 4966 -7342
rect 4883 -8301 4966 -7398
rect 43064 -7504 43400 -4872
rect 7504 -7672 43400 -7504
rect 3463 -8356 3880 -8344
rect 3463 -8412 3810 -8356
rect 3868 -8412 3880 -8356
rect 4883 -8357 4895 -8301
rect 4951 -8357 4966 -8301
rect 4883 -8361 4966 -8357
rect 3463 -8420 3880 -8412
rect 4013 -8413 4113 -8406
rect 3291 -9383 3367 -9363
rect 3291 -9439 3302 -9383
rect 3358 -9439 3367 -9383
rect 3291 -10143 3367 -9439
rect 3291 -10199 3302 -10143
rect 3358 -10199 3367 -10143
rect 3291 -10248 3367 -10199
rect 3463 -10138 3539 -8420
rect 4013 -8469 4034 -8413
rect 4091 -8469 4113 -8413
rect 4013 -8478 4113 -8469
rect 7558 -9299 7634 -7672
rect 9762 -7736 9844 -7728
rect 9762 -7792 9775 -7736
rect 9831 -7792 9844 -7736
rect 9762 -8302 9844 -7792
rect 3670 -9317 3776 -9299
rect 3670 -9373 3696 -9317
rect 3752 -9373 3776 -9317
rect 7558 -9352 7569 -9299
rect 7623 -9352 7634 -9299
rect 7558 -9365 7634 -9352
rect 8391 -8358 8749 -8349
rect 8391 -8411 8656 -8358
rect 8714 -8411 8749 -8358
rect 9762 -8358 9775 -8302
rect 9831 -8358 9844 -8302
rect 9762 -8361 9844 -8358
rect 8391 -8427 8749 -8411
rect 8854 -8411 8968 -8405
rect 3670 -9397 3776 -9373
rect 7591 -9450 8083 -9439
rect 7591 -9451 8019 -9450
rect 7591 -9504 7602 -9451
rect 7656 -9503 8019 -9451
rect 8073 -9503 8083 -9450
rect 7656 -9504 8083 -9503
rect 7591 -9515 8083 -9504
rect 7798 -9856 7874 -9515
rect 8391 -9735 8467 -8427
rect 8854 -8471 8878 -8411
rect 8942 -8471 8968 -8411
rect 8854 -8481 8968 -8471
rect 8529 -9307 8645 -9296
rect 8529 -9383 8566 -9307
rect 8627 -9383 8645 -9307
rect 12404 -9299 12480 -7672
rect 14570 -7733 14655 -7728
rect 14570 -7789 14584 -7733
rect 14640 -7789 14655 -7733
rect 14570 -8302 14655 -7789
rect 12404 -9352 12415 -9299
rect 12469 -9352 12480 -9299
rect 12404 -9365 12480 -9352
rect 13236 -8359 13588 -8349
rect 13236 -8411 13500 -8359
rect 13561 -8411 13588 -8359
rect 14570 -8358 14584 -8302
rect 14640 -8358 14655 -8302
rect 14570 -8361 14655 -8358
rect 13236 -8427 13588 -8411
rect 13705 -8413 13804 -8401
rect 8529 -9402 8645 -9383
rect 12437 -9450 12929 -9439
rect 12437 -9451 12865 -9450
rect 12437 -9504 12448 -9451
rect 12502 -9503 12865 -9451
rect 12919 -9503 12929 -9450
rect 12502 -9504 12929 -9503
rect 12437 -9515 12929 -9504
rect 8391 -9791 8401 -9735
rect 8457 -9791 8467 -9735
rect 8391 -9797 8467 -9791
rect 12644 -9856 12720 -9515
rect 13236 -9732 13313 -8427
rect 13705 -8469 13726 -8413
rect 13782 -8469 13804 -8413
rect 13705 -8478 13804 -8469
rect 13467 -9314 13579 -9296
rect 13467 -9373 13505 -9314
rect 13570 -9373 13579 -9314
rect 17250 -9299 17326 -7672
rect 19448 -7736 19531 -7728
rect 19448 -7792 19462 -7736
rect 19518 -7792 19531 -7736
rect 19448 -8301 19531 -7792
rect 17250 -9352 17261 -9299
rect 17315 -9352 17326 -9299
rect 17250 -9365 17326 -9352
rect 18078 -8357 18431 -8349
rect 18078 -8412 18347 -8357
rect 18407 -8412 18431 -8357
rect 19448 -8357 19460 -8301
rect 19516 -8357 19531 -8301
rect 19448 -8361 19531 -8357
rect 18078 -8427 18431 -8412
rect 18550 -8412 18647 -8398
rect 13467 -9399 13579 -9373
rect 17283 -9450 17775 -9439
rect 17283 -9451 17711 -9450
rect 17283 -9504 17294 -9451
rect 17348 -9503 17711 -9451
rect 17765 -9503 17775 -9450
rect 17348 -9504 17775 -9503
rect 17283 -9515 17775 -9504
rect 13236 -9788 13245 -9732
rect 13301 -9788 13313 -9732
rect 13236 -9796 13313 -9788
rect 17490 -9856 17566 -9515
rect 18078 -9734 18154 -8427
rect 18550 -8470 18571 -8412
rect 18629 -8470 18647 -8412
rect 18550 -8493 18647 -8470
rect 18226 -9317 18333 -9296
rect 18226 -9376 18252 -9317
rect 18318 -9376 18333 -9317
rect 22096 -9299 22172 -7672
rect 24259 -7737 24344 -7728
rect 24259 -7793 24273 -7737
rect 24329 -7793 24344 -7737
rect 24259 -8301 24344 -7793
rect 22096 -9352 22107 -9299
rect 22161 -9352 22172 -9299
rect 22096 -9365 22172 -9352
rect 22951 -8359 23274 -8349
rect 22951 -8411 23196 -8359
rect 23251 -8411 23274 -8359
rect 24259 -8357 24273 -8301
rect 24329 -8357 24344 -8301
rect 24259 -8361 24344 -8357
rect 22951 -8427 23274 -8411
rect 23405 -8406 23490 -8393
rect 18226 -9396 18333 -9376
rect 22129 -9450 22621 -9439
rect 22129 -9451 22557 -9450
rect 22129 -9504 22140 -9451
rect 22194 -9503 22557 -9451
rect 22611 -9503 22621 -9450
rect 22194 -9504 22621 -9503
rect 22129 -9515 22621 -9504
rect 18078 -9790 18088 -9734
rect 18144 -9790 18154 -9734
rect 18078 -9797 18154 -9790
rect 22336 -9856 22412 -9515
rect 22951 -9740 23027 -8427
rect 23405 -8471 23416 -8406
rect 23479 -8471 23490 -8406
rect 23405 -8481 23490 -8471
rect 23153 -9314 23265 -9295
rect 23153 -9373 23194 -9314
rect 23252 -9373 23265 -9314
rect 26942 -9299 27018 -7672
rect 29135 -7734 29216 -7728
rect 29135 -7790 29149 -7734
rect 29205 -7790 29216 -7734
rect 29135 -8302 29216 -7790
rect 26942 -9352 26953 -9299
rect 27007 -9352 27018 -9299
rect 26942 -9365 27018 -9352
rect 27768 -8357 28117 -8342
rect 27768 -8409 28042 -8357
rect 28097 -8409 28117 -8357
rect 29135 -8358 29148 -8302
rect 29204 -8358 29216 -8302
rect 29135 -8361 29216 -8358
rect 27768 -8420 28117 -8409
rect 28247 -8411 28343 -8401
rect 23153 -9397 23265 -9373
rect 26975 -9450 27467 -9439
rect 26975 -9451 27403 -9450
rect 26975 -9504 26986 -9451
rect 27040 -9503 27403 -9451
rect 27457 -9503 27467 -9450
rect 27040 -9504 27467 -9503
rect 26975 -9515 27467 -9504
rect 22951 -9796 22961 -9740
rect 23017 -9796 23027 -9740
rect 22951 -9800 23027 -9796
rect 27182 -9856 27258 -9515
rect 27768 -9737 27844 -8420
rect 28247 -8469 28262 -8411
rect 28323 -8469 28343 -8411
rect 28247 -8487 28343 -8469
rect 27968 -9317 28077 -9293
rect 27968 -9375 27993 -9317
rect 28053 -9375 28077 -9317
rect 31788 -9299 31864 -7672
rect 33979 -7734 34061 -7728
rect 33979 -7790 33993 -7734
rect 34049 -7790 34061 -7734
rect 33979 -8302 34061 -7790
rect 31788 -9352 31799 -9299
rect 31853 -9352 31864 -9299
rect 31788 -9365 31864 -9352
rect 32636 -8360 33001 -8352
rect 32636 -8413 32886 -8360
rect 32943 -8413 33001 -8360
rect 33979 -8358 33992 -8302
rect 34048 -8358 34061 -8302
rect 33979 -8361 34061 -8358
rect 32636 -8430 33001 -8413
rect 33093 -8413 33183 -8403
rect 27968 -9397 28077 -9375
rect 31821 -9450 32313 -9439
rect 31821 -9451 32249 -9450
rect 31821 -9504 31832 -9451
rect 31886 -9503 32249 -9451
rect 32303 -9503 32313 -9450
rect 31886 -9504 32313 -9503
rect 31821 -9515 32313 -9504
rect 27768 -9793 27778 -9737
rect 27834 -9793 27844 -9737
rect 27768 -9800 27844 -9793
rect 32028 -9856 32104 -9515
rect 32636 -9739 32712 -8430
rect 33093 -8471 33107 -8413
rect 33166 -8471 33183 -8413
rect 33093 -8484 33183 -8471
rect 36634 -9299 36710 -7672
rect 38823 -7738 38903 -7728
rect 38823 -7794 38833 -7738
rect 38889 -7794 38903 -7738
rect 38823 -8301 38903 -7794
rect 38823 -8357 38835 -8301
rect 38891 -8357 38903 -8301
rect 38823 -8361 38903 -8357
rect 32853 -9316 32946 -9300
rect 32853 -9374 32867 -9316
rect 32933 -9374 32946 -9316
rect 36634 -9352 36645 -9299
rect 36699 -9352 36710 -9299
rect 36634 -9365 36710 -9352
rect 37455 -8414 38027 -8404
rect 37455 -8467 37957 -8414
rect 38012 -8467 38027 -8414
rect 37455 -8480 38027 -8467
rect 32853 -9387 32946 -9374
rect 36667 -9450 37159 -9439
rect 36667 -9451 37095 -9450
rect 36667 -9504 36678 -9451
rect 36732 -9503 37095 -9451
rect 37149 -9503 37159 -9450
rect 36732 -9504 37159 -9503
rect 36667 -9515 37159 -9504
rect 32636 -9795 32646 -9739
rect 32702 -9795 32712 -9739
rect 32636 -9800 32712 -9795
rect 36874 -9856 36950 -9515
rect 37455 -9736 37531 -8480
rect 41480 -9299 41556 -7672
rect 37734 -9315 37811 -9303
rect 37734 -9371 37744 -9315
rect 37800 -9371 37811 -9315
rect 41480 -9352 41491 -9299
rect 41545 -9352 41556 -9299
rect 41480 -9365 41556 -9352
rect 37734 -9381 37811 -9371
rect 41513 -9450 42005 -9439
rect 41513 -9451 41941 -9450
rect 41513 -9504 41524 -9451
rect 41578 -9503 41941 -9451
rect 41995 -9503 42005 -9450
rect 41578 -9504 42005 -9503
rect 41513 -9515 42005 -9504
rect 37455 -9792 37465 -9736
rect 37521 -9792 37531 -9736
rect 37455 -9796 37531 -9792
rect 41720 -9856 41796 -9515
rect 7392 -9912 42828 -9856
rect 7392 -9968 42672 -9912
rect 42728 -9968 42828 -9912
rect 7392 -10024 42828 -9968
rect 3463 -10194 3473 -10138
rect 3529 -10194 3539 -10138
rect 3463 -10248 3539 -10194
rect 4883 -10144 4966 -10080
rect 4883 -10200 4896 -10144
rect 4952 -10200 4966 -10144
rect 4883 -11100 4966 -10200
rect 43064 -10304 43400 -7672
rect 7504 -10472 43400 -10304
rect 4883 -11156 4895 -11100
rect 4951 -11156 4966 -11100
rect 4883 -11161 4966 -11156
rect 4013 -11212 4108 -11207
rect 3460 -11236 3895 -11227
rect 3460 -11292 3811 -11236
rect 3867 -11292 3895 -11236
rect 4013 -11268 4035 -11212
rect 4091 -11268 4108 -11212
rect 4013 -11277 4108 -11268
rect 3460 -11305 3895 -11292
rect 3090 -11421 3161 -11374
rect 3090 -11445 3096 -11421
rect 2860 -11514 3096 -11445
rect 3157 -11514 3161 -11421
rect 2860 -11517 3161 -11514
rect 2860 -11876 2932 -11517
rect 3090 -11527 3161 -11517
rect 2860 -11959 2865 -11876
rect 2926 -11959 2932 -11876
rect 2860 -11977 2932 -11959
rect 3182 -12169 3283 -12153
rect 3182 -12225 3203 -12169
rect 3259 -12225 3283 -12169
rect 3182 -12715 3283 -12225
rect 3182 -12945 3284 -12715
rect 3182 -13001 3205 -12945
rect 3261 -13001 3284 -12945
rect 3182 -13048 3284 -13001
rect 3460 -12940 3536 -11305
rect 3665 -12107 3777 -12095
rect 3665 -12183 3688 -12107
rect 3758 -12183 3777 -12107
rect 7558 -12099 7634 -10472
rect 9762 -10534 9844 -10528
rect 9762 -10590 9776 -10534
rect 9832 -10590 9844 -10534
rect 9762 -11101 9844 -10590
rect 7558 -12152 7569 -12099
rect 7623 -12152 7634 -12099
rect 7558 -12165 7634 -12152
rect 8391 -11156 8725 -11149
rect 8391 -11212 8654 -11156
rect 8710 -11212 8725 -11156
rect 9762 -11157 9776 -11101
rect 9832 -11157 9844 -11101
rect 9762 -11161 9844 -11157
rect 8391 -11221 8725 -11212
rect 8855 -11212 8956 -11201
rect 3665 -12198 3777 -12183
rect 7591 -12250 8083 -12239
rect 7591 -12251 8019 -12250
rect 7591 -12304 7602 -12251
rect 7656 -12303 8019 -12251
rect 8073 -12303 8083 -12250
rect 7656 -12304 8083 -12303
rect 7591 -12315 8083 -12304
rect 7798 -12656 7874 -12315
rect 8391 -12533 8467 -11221
rect 8855 -11272 8874 -11212
rect 8938 -11272 8956 -11212
rect 8855 -11284 8956 -11272
rect 8523 -12114 8641 -12093
rect 8523 -12174 8559 -12114
rect 8617 -12174 8641 -12114
rect 12404 -12099 12480 -10472
rect 14570 -10535 14655 -10528
rect 14570 -10591 14584 -10535
rect 14640 -10591 14655 -10535
rect 14570 -11102 14655 -10591
rect 12404 -12152 12415 -12099
rect 12469 -12152 12480 -12099
rect 12404 -12165 12480 -12152
rect 13240 -11158 13575 -11150
rect 13240 -11210 13502 -11158
rect 13557 -11210 13575 -11158
rect 14570 -11158 14586 -11102
rect 14642 -11158 14655 -11102
rect 14570 -11161 14655 -11158
rect 13240 -11215 13575 -11210
rect 13707 -11212 13797 -11202
rect 8523 -12204 8641 -12174
rect 12437 -12250 12929 -12239
rect 12437 -12251 12865 -12250
rect 12437 -12304 12448 -12251
rect 12502 -12303 12865 -12251
rect 12919 -12303 12929 -12250
rect 12502 -12304 12929 -12303
rect 12437 -12315 12929 -12304
rect 8391 -12589 8401 -12533
rect 8457 -12589 8467 -12533
rect 8391 -12598 8467 -12589
rect 12644 -12656 12720 -12315
rect 13240 -12529 13316 -11215
rect 13707 -11269 13726 -11212
rect 13782 -11269 13797 -11212
rect 13707 -11284 13797 -11269
rect 13474 -12116 13574 -12096
rect 13474 -12173 13504 -12116
rect 13564 -12173 13574 -12116
rect 17250 -12099 17326 -10472
rect 19448 -10535 19531 -10528
rect 19448 -10591 19462 -10535
rect 19518 -10591 19531 -10535
rect 19448 -11099 19531 -10591
rect 17250 -12152 17261 -12099
rect 17315 -12152 17326 -12099
rect 17250 -12165 17326 -12152
rect 18082 -11155 18421 -11147
rect 18082 -11209 18347 -11155
rect 18404 -11209 18421 -11155
rect 19448 -11155 19461 -11099
rect 19517 -11155 19531 -11099
rect 19448 -11161 19531 -11155
rect 18082 -11220 18421 -11209
rect 18556 -11210 18647 -11195
rect 13474 -12192 13574 -12173
rect 17283 -12250 17775 -12239
rect 17283 -12251 17711 -12250
rect 17283 -12304 17294 -12251
rect 17348 -12303 17711 -12251
rect 17765 -12303 17775 -12250
rect 17348 -12304 17775 -12303
rect 17283 -12315 17775 -12304
rect 13240 -12585 13250 -12529
rect 13306 -12585 13316 -12529
rect 13240 -12596 13316 -12585
rect 17490 -12656 17566 -12315
rect 18082 -12533 18158 -11220
rect 18556 -11270 18571 -11210
rect 18630 -11270 18647 -11210
rect 18556 -11284 18647 -11270
rect 18221 -12118 18325 -12094
rect 18221 -12177 18249 -12118
rect 18313 -12177 18325 -12118
rect 22096 -12099 22172 -10472
rect 24259 -10534 24344 -10528
rect 24259 -10590 24274 -10534
rect 24330 -10590 24344 -10534
rect 24259 -11100 24344 -10590
rect 22096 -12152 22107 -12099
rect 22161 -12152 22172 -12099
rect 22096 -12165 22172 -12152
rect 22922 -11156 23265 -11150
rect 22922 -11208 23194 -11156
rect 23253 -11208 23265 -11156
rect 24259 -11156 24274 -11100
rect 24330 -11156 24344 -11100
rect 24259 -11161 24344 -11156
rect 22922 -11213 23265 -11208
rect 23405 -11210 23490 -11197
rect 18221 -12198 18325 -12177
rect 22129 -12250 22621 -12239
rect 22129 -12251 22557 -12250
rect 22129 -12304 22140 -12251
rect 22194 -12303 22557 -12251
rect 22611 -12303 22621 -12250
rect 22194 -12304 22621 -12303
rect 22129 -12315 22621 -12304
rect 18082 -12589 18092 -12533
rect 18148 -12589 18158 -12533
rect 18082 -12597 18158 -12589
rect 22336 -12656 22412 -12315
rect 22922 -12537 22998 -11213
rect 23405 -11270 23417 -11210
rect 23480 -11270 23490 -11210
rect 23405 -11283 23490 -11270
rect 23150 -12113 23268 -12095
rect 23150 -12176 23190 -12113
rect 23255 -12176 23268 -12113
rect 26942 -12099 27018 -10472
rect 29135 -10533 29216 -10528
rect 29135 -10589 29147 -10533
rect 29203 -10589 29216 -10533
rect 29135 -11100 29216 -10589
rect 26942 -12152 26953 -12099
rect 27007 -12152 27018 -12099
rect 26942 -12165 27018 -12152
rect 27766 -11158 28122 -11149
rect 27766 -11212 28039 -11158
rect 28098 -11212 28122 -11158
rect 29135 -11156 29148 -11100
rect 29204 -11156 29216 -11100
rect 29135 -11161 29216 -11156
rect 27766 -11222 28122 -11212
rect 28248 -11212 28335 -11204
rect 23150 -12194 23268 -12176
rect 26975 -12250 27467 -12239
rect 26975 -12251 27403 -12250
rect 26975 -12304 26986 -12251
rect 27040 -12303 27403 -12251
rect 27457 -12303 27467 -12250
rect 27040 -12304 27467 -12303
rect 26975 -12315 27467 -12304
rect 22922 -12593 22932 -12537
rect 22988 -12593 22998 -12537
rect 22922 -12600 22998 -12593
rect 27182 -12656 27258 -12315
rect 27766 -12533 27842 -11222
rect 28248 -11268 28264 -11212
rect 28320 -11268 28335 -11212
rect 28248 -11278 28335 -11268
rect 31788 -12099 31864 -10472
rect 33979 -10536 34061 -10528
rect 33979 -10592 33992 -10536
rect 34048 -10592 34061 -10536
rect 33979 -11099 34061 -10592
rect 27977 -12117 28074 -12100
rect 27977 -12175 27998 -12117
rect 28058 -12175 28074 -12117
rect 31788 -12152 31799 -12099
rect 31853 -12152 31864 -12099
rect 31788 -12165 31864 -12152
rect 32638 -11156 32959 -11150
rect 32638 -11211 32888 -11156
rect 32947 -11211 32959 -11156
rect 33979 -11155 33993 -11099
rect 34049 -11155 34061 -11099
rect 33979 -11161 34061 -11155
rect 32638 -11221 32959 -11211
rect 33095 -11212 33179 -11203
rect 27977 -12195 28074 -12175
rect 31821 -12250 32313 -12239
rect 31821 -12251 32249 -12250
rect 31821 -12304 31832 -12251
rect 31886 -12303 32249 -12251
rect 32303 -12303 32313 -12250
rect 31886 -12304 32313 -12303
rect 31821 -12315 32313 -12304
rect 27766 -12589 27776 -12533
rect 27832 -12589 27842 -12533
rect 27766 -12598 27842 -12589
rect 32028 -12656 32104 -12315
rect 32638 -12536 32714 -11221
rect 33095 -11268 33111 -11212
rect 33167 -11268 33179 -11212
rect 33095 -11279 33179 -11268
rect 36634 -12099 36710 -10472
rect 38823 -10534 38903 -10528
rect 38823 -10590 38836 -10534
rect 38892 -10590 38903 -10534
rect 38823 -11100 38903 -10590
rect 38823 -11156 38835 -11100
rect 38891 -11156 38903 -11100
rect 38823 -11161 38903 -11156
rect 32865 -12116 32956 -12100
rect 32865 -12173 32888 -12116
rect 32944 -12173 32956 -12116
rect 36634 -12152 36645 -12099
rect 36699 -12152 36710 -12099
rect 36634 -12165 36710 -12152
rect 37456 -11212 38024 -11203
rect 37456 -11268 37957 -11212
rect 38013 -11268 38024 -11212
rect 37456 -11279 38024 -11268
rect 32865 -12190 32956 -12173
rect 36667 -12250 37159 -12239
rect 36667 -12251 37095 -12250
rect 36667 -12304 36678 -12251
rect 36732 -12303 37095 -12251
rect 37149 -12303 37159 -12250
rect 36732 -12304 37159 -12303
rect 36667 -12315 37159 -12304
rect 32638 -12592 32648 -12536
rect 32704 -12592 32714 -12536
rect 32638 -12599 32714 -12592
rect 36874 -12656 36950 -12315
rect 37456 -12534 37532 -11279
rect 41480 -12099 41556 -10472
rect 37731 -12114 37811 -12103
rect 37731 -12170 37744 -12114
rect 37800 -12170 37811 -12114
rect 41480 -12152 41491 -12099
rect 41545 -12152 41556 -12099
rect 41480 -12165 41556 -12152
rect 37731 -12182 37811 -12170
rect 41513 -12250 42005 -12239
rect 41513 -12251 41941 -12250
rect 41513 -12304 41524 -12251
rect 41578 -12303 41941 -12251
rect 41995 -12303 42005 -12250
rect 41578 -12304 42005 -12303
rect 41513 -12315 42005 -12304
rect 37456 -12590 37466 -12534
rect 37522 -12590 37532 -12534
rect 37456 -12597 37532 -12590
rect 41720 -12656 41796 -12315
rect 7392 -12712 42841 -12656
rect 7392 -12768 42672 -12712
rect 42728 -12768 42841 -12712
rect 7392 -12824 42841 -12768
rect 3460 -12996 3469 -12940
rect 3525 -12996 3536 -12940
rect 3460 -13048 3536 -12996
rect 4883 -12940 4966 -12880
rect 4883 -12996 4895 -12940
rect 4951 -12996 4966 -12940
rect 4883 -13902 4966 -12996
rect 43064 -13104 43400 -10472
rect 7504 -13272 43400 -13104
rect 4883 -13958 4895 -13902
rect 4951 -13958 4966 -13902
rect 4883 -13961 4966 -13958
rect 4015 -14013 4108 -14001
rect 3461 -14035 3920 -14028
rect 3461 -14088 3808 -14035
rect 3871 -14088 3920 -14035
rect 4015 -14070 4035 -14013
rect 4092 -14070 4108 -14013
rect 4015 -14078 4108 -14070
rect 3461 -14105 3920 -14088
rect 3167 -14907 3269 -14893
rect 3167 -14963 3187 -14907
rect 3243 -14963 3269 -14907
rect 3167 -15738 3269 -14963
rect 3167 -15794 3191 -15738
rect 3247 -15794 3269 -15738
rect 3167 -15848 3269 -15794
rect 3461 -15746 3537 -14105
rect 3656 -14907 3771 -14898
rect 3656 -14983 3681 -14907
rect 3746 -14983 3771 -14907
rect 7558 -14899 7634 -13272
rect 9762 -13340 9844 -13328
rect 9762 -13396 9774 -13340
rect 9830 -13396 9844 -13340
rect 9762 -13901 9844 -13396
rect 7558 -14952 7569 -14899
rect 7623 -14952 7634 -14899
rect 7558 -14965 7634 -14952
rect 8392 -13957 8734 -13948
rect 8392 -14012 8657 -13957
rect 8712 -14012 8734 -13957
rect 9762 -13957 9775 -13901
rect 9831 -13957 9844 -13901
rect 9762 -13961 9844 -13957
rect 8392 -14020 8734 -14012
rect 8850 -14011 8968 -13998
rect 3656 -14995 3771 -14983
rect 7591 -15050 8083 -15039
rect 7591 -15051 8019 -15050
rect 7591 -15104 7602 -15051
rect 7656 -15103 8019 -15051
rect 8073 -15103 8083 -15050
rect 7656 -15104 8083 -15103
rect 7591 -15115 8083 -15104
rect 7798 -15456 7874 -15115
rect 8392 -15337 8468 -14020
rect 8850 -14069 8879 -14011
rect 8939 -14069 8968 -14011
rect 8850 -14080 8968 -14069
rect 8539 -14917 8649 -14896
rect 8539 -14973 8578 -14917
rect 8636 -14973 8649 -14917
rect 12404 -14899 12480 -13272
rect 14570 -13335 14655 -13328
rect 14570 -13391 14583 -13335
rect 14639 -13391 14655 -13335
rect 14570 -13902 14655 -13391
rect 12404 -14952 12415 -14899
rect 12469 -14952 12480 -14899
rect 12404 -14965 12480 -14952
rect 13238 -13956 13586 -13949
rect 13238 -14010 13504 -13956
rect 13559 -14010 13586 -13956
rect 14570 -13958 14585 -13902
rect 14641 -13958 14655 -13902
rect 14570 -13961 14655 -13958
rect 13238 -14025 13586 -14010
rect 13707 -14012 13799 -14005
rect 8539 -14997 8649 -14973
rect 12437 -15050 12929 -15039
rect 12437 -15051 12865 -15050
rect 12437 -15104 12448 -15051
rect 12502 -15103 12865 -15051
rect 12919 -15103 12929 -15050
rect 12502 -15104 12929 -15103
rect 12437 -15115 12929 -15104
rect 8392 -15393 8402 -15337
rect 8458 -15393 8468 -15337
rect 8392 -15400 8468 -15393
rect 12644 -15456 12720 -15115
rect 13238 -15339 13314 -14025
rect 13707 -14069 13725 -14012
rect 13784 -14069 13799 -14012
rect 13707 -14079 13799 -14069
rect 13474 -14916 13578 -14897
rect 13474 -14973 13509 -14916
rect 13568 -14973 13578 -14916
rect 17250 -14899 17326 -13272
rect 19448 -13333 19531 -13328
rect 19448 -13389 19461 -13333
rect 19517 -13389 19531 -13333
rect 19448 -13900 19531 -13389
rect 17250 -14952 17261 -14899
rect 17315 -14952 17326 -14899
rect 17250 -14965 17326 -14952
rect 18081 -13955 18430 -13946
rect 18081 -14011 18348 -13955
rect 18406 -14011 18430 -13955
rect 19448 -13956 19462 -13900
rect 19518 -13956 19531 -13900
rect 19448 -13961 19531 -13956
rect 18081 -14024 18430 -14011
rect 18551 -14011 18649 -13996
rect 13474 -14991 13578 -14973
rect 17283 -15050 17775 -15039
rect 17283 -15051 17711 -15050
rect 17283 -15104 17294 -15051
rect 17348 -15103 17711 -15051
rect 17765 -15103 17775 -15050
rect 17348 -15104 17775 -15103
rect 17283 -15115 17775 -15104
rect 13238 -15395 13248 -15339
rect 13304 -15395 13314 -15339
rect 13238 -15400 13314 -15395
rect 17490 -15456 17566 -15115
rect 18081 -15335 18157 -14024
rect 18551 -14068 18572 -14011
rect 18630 -14068 18649 -14011
rect 18551 -14088 18649 -14068
rect 18227 -14917 18340 -14891
rect 18227 -14979 18252 -14917
rect 18316 -14979 18340 -14917
rect 22096 -14899 22172 -13272
rect 24259 -13334 24344 -13328
rect 24259 -13390 24275 -13334
rect 24331 -13390 24344 -13334
rect 24259 -13901 24344 -13390
rect 22096 -14952 22107 -14899
rect 22161 -14952 22172 -14899
rect 22096 -14965 22172 -14952
rect 22950 -13957 23271 -13946
rect 22950 -14011 23196 -13957
rect 23255 -14011 23271 -13957
rect 24259 -13957 24274 -13901
rect 24330 -13957 24344 -13901
rect 24259 -13961 24344 -13957
rect 22950 -14020 23271 -14011
rect 23405 -14013 23488 -14001
rect 18227 -15005 18340 -14979
rect 22129 -15050 22621 -15039
rect 22129 -15051 22557 -15050
rect 22129 -15104 22140 -15051
rect 22194 -15103 22557 -15051
rect 22611 -15103 22621 -15050
rect 22194 -15104 22621 -15103
rect 22129 -15115 22621 -15104
rect 18081 -15391 18091 -15335
rect 18147 -15391 18157 -15335
rect 18081 -15397 18157 -15391
rect 22336 -15456 22412 -15115
rect 22950 -15335 23026 -14020
rect 23405 -14070 23417 -14013
rect 23477 -14070 23488 -14013
rect 23405 -14080 23488 -14070
rect 23147 -14909 23265 -14892
rect 23147 -14974 23191 -14909
rect 23254 -14974 23265 -14909
rect 26942 -14899 27018 -13272
rect 29135 -13332 29216 -13328
rect 29135 -13388 29148 -13332
rect 29204 -13388 29216 -13332
rect 29135 -13900 29216 -13388
rect 27765 -13950 28122 -13942
rect 27765 -14012 28039 -13950
rect 28099 -14012 28122 -13950
rect 29135 -13956 29147 -13900
rect 29203 -13956 29216 -13900
rect 29135 -13961 29216 -13956
rect 27765 -14023 28122 -14012
rect 28250 -14012 28333 -14003
rect 26942 -14952 26953 -14899
rect 27007 -14952 27018 -14899
rect 26942 -14965 27018 -14952
rect 23147 -14996 23265 -14974
rect 26975 -15050 27467 -15039
rect 26975 -15051 27403 -15050
rect 26975 -15104 26986 -15051
rect 27040 -15103 27403 -15051
rect 27457 -15103 27467 -15050
rect 27040 -15104 27467 -15103
rect 26975 -15115 27467 -15104
rect 22950 -15391 22960 -15335
rect 23016 -15391 23026 -15335
rect 22950 -15396 23026 -15391
rect 27182 -15456 27258 -15115
rect 27767 -15335 27843 -14023
rect 28250 -14068 28263 -14012
rect 28321 -14068 28333 -14012
rect 28250 -14076 28333 -14068
rect 31788 -14899 31864 -13272
rect 33979 -13335 34061 -13328
rect 33979 -13391 33993 -13335
rect 34049 -13391 34061 -13335
rect 33979 -13900 34061 -13391
rect 27979 -14916 28076 -14899
rect 27979 -14972 27997 -14916
rect 28062 -14972 28076 -14916
rect 31788 -14952 31799 -14899
rect 31853 -14952 31864 -14899
rect 31788 -14965 31864 -14952
rect 32638 -13955 32967 -13948
rect 32638 -14014 32885 -13955
rect 32947 -14014 32967 -13955
rect 33979 -13956 33991 -13900
rect 34047 -13956 34061 -13900
rect 33979 -13961 34061 -13956
rect 32638 -14023 32967 -14014
rect 33095 -14012 33178 -14005
rect 27979 -14989 28076 -14972
rect 31821 -15050 32313 -15039
rect 31821 -15051 32249 -15050
rect 31821 -15104 31832 -15051
rect 31886 -15103 32249 -15051
rect 32303 -15103 32313 -15050
rect 31886 -15104 32313 -15103
rect 31821 -15115 32313 -15104
rect 27767 -15391 27777 -15335
rect 27833 -15391 27843 -15335
rect 27767 -15396 27843 -15391
rect 32028 -15456 32104 -15115
rect 32638 -15332 32714 -14023
rect 33095 -14069 33110 -14012
rect 33166 -14069 33178 -14012
rect 33095 -14078 33178 -14069
rect 36634 -14899 36710 -13272
rect 38823 -13335 38903 -13328
rect 38823 -13391 38837 -13335
rect 38893 -13391 38903 -13335
rect 38823 -13901 38903 -13391
rect 38823 -13957 38835 -13901
rect 38891 -13957 38903 -13901
rect 38823 -13961 38903 -13957
rect 32845 -14916 32949 -14904
rect 32845 -14974 32866 -14916
rect 32938 -14974 32949 -14916
rect 36634 -14952 36645 -14899
rect 36699 -14952 36710 -14899
rect 36634 -14965 36710 -14952
rect 37454 -14013 38025 -14002
rect 37454 -14067 37957 -14013
rect 38013 -14067 38025 -14013
rect 37454 -14078 38025 -14067
rect 32845 -14989 32949 -14974
rect 36667 -15050 37159 -15039
rect 36667 -15051 37095 -15050
rect 36667 -15104 36678 -15051
rect 36732 -15103 37095 -15051
rect 37149 -15103 37159 -15050
rect 36732 -15104 37159 -15103
rect 36667 -15115 37159 -15104
rect 32638 -15388 32648 -15332
rect 32704 -15388 32714 -15332
rect 32638 -15396 32714 -15388
rect 36874 -15456 36950 -15115
rect 37454 -15331 37530 -14078
rect 41480 -14899 41556 -13272
rect 37733 -14914 37812 -14903
rect 37733 -14970 37744 -14914
rect 37800 -14970 37812 -14914
rect 41480 -14952 41491 -14899
rect 41545 -14952 41556 -14899
rect 41480 -14965 41556 -14952
rect 37733 -14981 37812 -14970
rect 41513 -15050 42005 -15039
rect 41513 -15051 41941 -15050
rect 41513 -15104 41524 -15051
rect 41578 -15103 41941 -15051
rect 41995 -15103 42005 -15050
rect 41578 -15104 42005 -15103
rect 41513 -15115 42005 -15104
rect 37454 -15387 37464 -15331
rect 37520 -15387 37530 -15331
rect 37454 -15396 37530 -15387
rect 41720 -15456 41796 -15115
rect 7392 -15512 42868 -15456
rect 7392 -15568 42672 -15512
rect 42728 -15568 42868 -15512
rect 7392 -15624 42868 -15568
rect 3461 -15802 3471 -15746
rect 3527 -15802 3537 -15746
rect 3461 -15848 3537 -15802
rect 4883 -15740 4966 -15680
rect 4883 -15796 4898 -15740
rect 4954 -15796 4966 -15740
rect 4883 -16700 4966 -15796
rect 43064 -15904 43400 -13272
rect 7504 -16072 43400 -15904
rect 4883 -16756 4897 -16700
rect 4953 -16756 4966 -16700
rect 4883 -16761 4966 -16756
rect 3174 -16806 3256 -16779
rect 3174 -16883 3181 -16806
rect 3251 -16883 3256 -16806
rect 4018 -16812 4107 -16806
rect 3174 -16910 3256 -16883
rect 3462 -16829 3538 -16828
rect 3462 -16835 3917 -16829
rect 3462 -16891 3809 -16835
rect 3865 -16891 3917 -16835
rect 4018 -16868 4034 -16812
rect 4090 -16868 4107 -16812
rect 4018 -16876 4107 -16868
rect 3462 -16905 3917 -16891
rect 3180 -17099 3252 -16910
rect 2844 -17171 3256 -17099
rect 2844 -17716 2916 -17171
rect 2844 -17778 2850 -17716
rect 2911 -17778 2916 -17716
rect 2844 -17790 2916 -17778
rect 3462 -18513 3538 -16905
rect 3664 -17707 3776 -17696
rect 3664 -17783 3692 -17707
rect 3760 -17783 3776 -17707
rect 7558 -17699 7634 -16072
rect 9762 -16140 9844 -16128
rect 9762 -16196 9774 -16140
rect 9830 -16196 9844 -16140
rect 9762 -16700 9844 -16196
rect 7558 -17752 7569 -17699
rect 7623 -17752 7634 -17699
rect 7558 -17765 7634 -17752
rect 8390 -16757 8726 -16751
rect 8390 -16811 8654 -16757
rect 8713 -16811 8726 -16757
rect 9762 -16756 9775 -16700
rect 9831 -16756 9844 -16700
rect 9762 -16761 9844 -16756
rect 8390 -16816 8726 -16811
rect 8857 -16812 8959 -16805
rect 3664 -17796 3776 -17783
rect 7591 -17850 8083 -17839
rect 7591 -17851 8019 -17850
rect 7591 -17904 7602 -17851
rect 7656 -17903 8019 -17851
rect 8073 -17903 8083 -17850
rect 7656 -17904 8083 -17903
rect 7591 -17915 8083 -17904
rect 7798 -18256 7874 -17915
rect 8390 -18137 8466 -16816
rect 8857 -16870 8879 -16812
rect 8938 -16870 8959 -16812
rect 8857 -16879 8959 -16870
rect 8538 -17717 8646 -17693
rect 8538 -17775 8570 -17717
rect 8630 -17775 8646 -17717
rect 12404 -17699 12480 -16072
rect 14570 -16137 14655 -16128
rect 14570 -16193 14584 -16137
rect 14640 -16193 14655 -16137
rect 14570 -16701 14655 -16193
rect 12404 -17752 12415 -17699
rect 12469 -17752 12480 -17699
rect 12404 -17765 12480 -17752
rect 13252 -16754 13573 -16751
rect 13252 -16811 13501 -16754
rect 13560 -16811 13573 -16754
rect 14570 -16757 14585 -16701
rect 14641 -16757 14655 -16701
rect 14570 -16761 14655 -16757
rect 13252 -16814 13573 -16811
rect 13710 -16812 13795 -16806
rect 8538 -17798 8646 -17775
rect 12437 -17850 12929 -17839
rect 12437 -17851 12865 -17850
rect 12437 -17904 12448 -17851
rect 12502 -17903 12865 -17851
rect 12919 -17903 12929 -17850
rect 12502 -17904 12929 -17903
rect 12437 -17915 12929 -17904
rect 8390 -18193 8400 -18137
rect 8456 -18193 8466 -18137
rect 8390 -18200 8466 -18193
rect 12644 -18256 12720 -17915
rect 13252 -18140 13328 -16814
rect 13710 -16869 13726 -16812
rect 13785 -16869 13795 -16812
rect 13710 -16881 13795 -16869
rect 17250 -17699 17326 -16072
rect 19448 -16135 19531 -16128
rect 19448 -16191 19463 -16135
rect 19519 -16191 19531 -16135
rect 19448 -16701 19531 -16191
rect 13483 -17715 13572 -17699
rect 13483 -17771 13505 -17715
rect 13561 -17771 13572 -17715
rect 17250 -17752 17261 -17699
rect 17315 -17752 17326 -17699
rect 17250 -17765 17326 -17752
rect 18080 -16758 18434 -16752
rect 18080 -16815 18346 -16758
rect 18407 -16815 18434 -16758
rect 19448 -16757 19462 -16701
rect 19518 -16757 19531 -16701
rect 19448 -16761 19531 -16757
rect 18080 -16821 18434 -16815
rect 18558 -16810 18643 -16799
rect 13483 -17793 13572 -17771
rect 17283 -17850 17775 -17839
rect 17283 -17851 17711 -17850
rect 17283 -17904 17294 -17851
rect 17348 -17903 17711 -17851
rect 17765 -17903 17775 -17850
rect 17348 -17904 17775 -17903
rect 17283 -17915 17775 -17904
rect 13252 -18196 13262 -18140
rect 13318 -18196 13328 -18140
rect 13252 -18200 13328 -18196
rect 17490 -18256 17566 -17915
rect 18080 -18134 18156 -16821
rect 18558 -16869 18572 -16810
rect 18630 -16869 18643 -16810
rect 18558 -16884 18643 -16869
rect 18221 -17715 18335 -17695
rect 18221 -17776 18250 -17715
rect 18318 -17776 18335 -17715
rect 22096 -17699 22172 -16072
rect 24259 -16142 24344 -16128
rect 24259 -16198 24273 -16142
rect 24329 -16198 24344 -16142
rect 24259 -16702 24344 -16198
rect 22096 -17752 22107 -17699
rect 22161 -17752 22172 -17699
rect 22096 -17765 22172 -17752
rect 22946 -16757 23264 -16748
rect 22946 -16811 23194 -16757
rect 23252 -16811 23264 -16757
rect 24259 -16758 24274 -16702
rect 24330 -16758 24344 -16702
rect 24259 -16761 24344 -16758
rect 22946 -16815 23264 -16811
rect 23406 -16811 23491 -16801
rect 18221 -17796 18335 -17776
rect 22129 -17850 22621 -17839
rect 22129 -17851 22557 -17850
rect 22129 -17904 22140 -17851
rect 22194 -17903 22557 -17851
rect 22611 -17903 22621 -17850
rect 22194 -17904 22621 -17903
rect 22129 -17915 22621 -17904
rect 18080 -18190 18090 -18134
rect 18146 -18190 18156 -18134
rect 18080 -18195 18156 -18190
rect 22336 -18256 22412 -17915
rect 22946 -18134 23022 -16815
rect 23406 -16870 23415 -16811
rect 23478 -16870 23491 -16811
rect 23406 -16880 23491 -16870
rect 23153 -17712 23267 -17694
rect 23153 -17778 23191 -17712
rect 23251 -17778 23267 -17712
rect 26942 -17699 27018 -16072
rect 29135 -16134 29216 -16128
rect 29135 -16190 29148 -16134
rect 29204 -16190 29216 -16134
rect 29135 -16702 29216 -16190
rect 26942 -17752 26953 -17699
rect 27007 -17752 27018 -17699
rect 26942 -17765 27018 -17752
rect 27769 -16754 28115 -16749
rect 27769 -16811 28037 -16754
rect 28101 -16811 28115 -16754
rect 29135 -16758 29148 -16702
rect 29204 -16758 29216 -16702
rect 29135 -16761 29216 -16758
rect 27769 -16823 28115 -16811
rect 28249 -16811 28334 -16804
rect 23153 -17798 23267 -17778
rect 26975 -17850 27467 -17839
rect 26975 -17851 27403 -17850
rect 26975 -17904 26986 -17851
rect 27040 -17903 27403 -17851
rect 27457 -17903 27467 -17850
rect 27040 -17904 27467 -17903
rect 26975 -17915 27467 -17904
rect 22946 -18190 22956 -18134
rect 23012 -18190 23022 -18134
rect 22946 -18197 23022 -18190
rect 27182 -18256 27258 -17915
rect 27769 -18136 27845 -16823
rect 28249 -16867 28265 -16811
rect 28323 -16867 28334 -16811
rect 28249 -16875 28334 -16867
rect 27983 -17712 28077 -17698
rect 27983 -17769 27999 -17712
rect 28060 -17769 28077 -17712
rect 31788 -17699 31864 -16072
rect 33979 -16134 34061 -16128
rect 33979 -16190 33993 -16134
rect 34049 -16190 34061 -16134
rect 33979 -16700 34061 -16190
rect 31788 -17752 31799 -17699
rect 31853 -17752 31864 -17699
rect 31788 -17765 31864 -17752
rect 32636 -16755 32966 -16747
rect 32636 -16811 32884 -16755
rect 32943 -16811 32966 -16755
rect 33979 -16756 33993 -16700
rect 34049 -16756 34061 -16700
rect 33979 -16761 34061 -16756
rect 32636 -16819 32966 -16811
rect 33096 -16813 33184 -16801
rect 27983 -17787 28077 -17769
rect 31821 -17850 32313 -17839
rect 31821 -17851 32249 -17850
rect 31821 -17904 31832 -17851
rect 31886 -17903 32249 -17851
rect 32303 -17903 32313 -17850
rect 31886 -17904 32313 -17903
rect 31821 -17915 32313 -17904
rect 27769 -18192 27779 -18136
rect 27835 -18192 27845 -18136
rect 27769 -18198 27845 -18192
rect 32028 -18256 32104 -17915
rect 32636 -18138 32712 -16819
rect 33096 -16870 33109 -16813
rect 33167 -16870 33184 -16813
rect 33096 -16878 33184 -16870
rect 36634 -17699 36710 -16072
rect 38823 -16135 38903 -16128
rect 38823 -16191 38835 -16135
rect 38891 -16191 38903 -16135
rect 38823 -16701 38903 -16191
rect 38823 -16757 38835 -16701
rect 38891 -16757 38903 -16701
rect 38823 -16761 38903 -16757
rect 32850 -17715 32945 -17702
rect 32850 -17775 32868 -17715
rect 32935 -17775 32945 -17715
rect 36634 -17752 36645 -17699
rect 36699 -17752 36710 -17699
rect 36634 -17765 36710 -17752
rect 37456 -16812 38026 -16798
rect 37456 -16870 37952 -16812
rect 38016 -16870 38026 -16812
rect 37456 -16880 38026 -16870
rect 32850 -17791 32945 -17775
rect 36667 -17850 37159 -17839
rect 36667 -17851 37095 -17850
rect 36667 -17904 36678 -17851
rect 36732 -17903 37095 -17851
rect 37149 -17903 37159 -17850
rect 36732 -17904 37159 -17903
rect 36667 -17915 37159 -17904
rect 32636 -18194 32646 -18138
rect 32702 -18194 32712 -18138
rect 32636 -18199 32712 -18194
rect 36874 -18256 36950 -17915
rect 37456 -18197 37532 -16880
rect 41480 -17699 41556 -16072
rect 37735 -17716 37813 -17703
rect 37735 -17772 37744 -17716
rect 37800 -17772 37813 -17716
rect 41480 -17752 41491 -17699
rect 41545 -17752 41556 -17699
rect 41480 -17765 41556 -17752
rect 37735 -17783 37813 -17772
rect 41513 -17850 42005 -17839
rect 41513 -17851 41941 -17850
rect 41513 -17904 41524 -17851
rect 41578 -17903 41941 -17851
rect 41995 -17903 42005 -17850
rect 41578 -17904 42005 -17903
rect 41513 -17915 42005 -17904
rect 41720 -18256 41796 -17915
rect 7392 -18312 42841 -18256
rect 7392 -18368 42672 -18312
rect 42728 -18368 42841 -18312
rect 7392 -18424 42841 -18368
rect 3462 -18569 3471 -18513
rect 3527 -18569 3538 -18513
rect 3462 -18648 3538 -18569
rect 43064 -18704 43400 -16072
rect 7504 -18872 43400 -18704
rect 4872 -19499 4984 -19497
rect 4872 -19555 4893 -19499
rect 4956 -19555 4984 -19499
rect 4872 -19561 4984 -19555
rect 4018 -19613 4107 -19608
rect 4018 -19669 4034 -19613
rect 4091 -19669 4107 -19613
rect 4018 -19678 4107 -19669
rect 3664 -20507 3772 -20496
rect 3664 -20583 3696 -20507
rect 3752 -20583 3772 -20507
rect 7558 -20499 7634 -18872
rect 9744 -19498 9856 -19497
rect 9744 -19554 9772 -19498
rect 9834 -19554 9856 -19498
rect 9744 -19561 9856 -19554
rect 8862 -19612 8956 -19603
rect 8862 -19668 8881 -19612
rect 8939 -19668 8956 -19612
rect 8862 -19678 8956 -19668
rect 7558 -20552 7569 -20499
rect 7623 -20552 7634 -20499
rect 7558 -20565 7634 -20552
rect 8532 -20514 8651 -20494
rect 3664 -20596 3772 -20583
rect 8532 -20573 8563 -20514
rect 8625 -20573 8651 -20514
rect 12404 -20499 12480 -18872
rect 14560 -19501 14672 -19497
rect 14560 -19557 14580 -19501
rect 14645 -19557 14672 -19501
rect 14560 -19561 14672 -19557
rect 13713 -19612 13794 -19602
rect 13713 -19668 13727 -19612
rect 13784 -19668 13794 -19612
rect 13713 -19676 13794 -19668
rect 12404 -20552 12415 -20499
rect 12469 -20552 12480 -20499
rect 17250 -20499 17326 -18872
rect 19432 -19502 19544 -19497
rect 19432 -19558 19458 -19502
rect 19521 -19558 19544 -19502
rect 19432 -19561 19544 -19558
rect 18555 -19613 18649 -19595
rect 18555 -19669 18573 -19613
rect 18630 -19669 18649 -19613
rect 18555 -19683 18649 -19669
rect 12404 -20565 12480 -20552
rect 13484 -20515 13581 -20501
rect 8532 -20601 8651 -20573
rect 13484 -20571 13513 -20515
rect 13571 -20571 13581 -20515
rect 17250 -20552 17261 -20499
rect 17315 -20552 17326 -20499
rect 17250 -20565 17326 -20552
rect 18223 -20518 18334 -20497
rect 13484 -20589 13581 -20571
rect 18223 -20580 18251 -20518
rect 18315 -20580 18334 -20518
rect 22096 -20499 22172 -18872
rect 24248 -19499 24360 -19497
rect 24248 -19556 24269 -19499
rect 24334 -19556 24360 -19499
rect 24248 -19561 24360 -19556
rect 23404 -19612 23485 -19605
rect 23404 -19669 23417 -19612
rect 23476 -19669 23485 -19612
rect 23404 -19679 23485 -19669
rect 22096 -20552 22107 -20499
rect 22161 -20552 22172 -20499
rect 22096 -20565 22172 -20552
rect 23162 -20514 23270 -20496
rect 18223 -20598 18334 -20580
rect 23162 -20577 23193 -20514
rect 23253 -20577 23270 -20514
rect 26942 -20499 27018 -18872
rect 29120 -19502 29232 -19497
rect 29120 -19558 29145 -19502
rect 29206 -19558 29232 -19502
rect 29120 -19561 29232 -19558
rect 28246 -19612 28338 -19599
rect 28246 -19669 28262 -19612
rect 28319 -19669 28338 -19612
rect 28246 -19681 28338 -19669
rect 26942 -20552 26953 -20499
rect 27007 -20552 27018 -20499
rect 26942 -20565 27018 -20552
rect 27983 -20517 28072 -20496
rect 23162 -20597 23270 -20577
rect 27983 -20574 27998 -20517
rect 28059 -20574 28072 -20517
rect 31788 -20499 31864 -18872
rect 33963 -19501 34077 -19497
rect 33963 -19557 33989 -19501
rect 34051 -19557 34077 -19501
rect 33963 -19561 34077 -19557
rect 33090 -19611 33189 -19600
rect 33090 -19670 33108 -19611
rect 33170 -19670 33189 -19611
rect 33090 -19685 33189 -19670
rect 31788 -20552 31799 -20499
rect 31853 -20552 31864 -20499
rect 36634 -20499 36710 -18872
rect 38744 -18873 38996 -18872
rect 43064 -19219 43400 -18872
rect 31788 -20565 31864 -20552
rect 32859 -20517 32943 -20503
rect 27983 -20587 28072 -20574
rect 32859 -20574 32869 -20517
rect 32932 -20574 32943 -20517
rect 36634 -20552 36645 -20499
rect 36699 -20552 36710 -20499
rect 36634 -20565 36710 -20552
rect 32859 -20586 32943 -20574
rect 7591 -20650 8083 -20639
rect 7591 -20651 8019 -20650
rect 7591 -20704 7602 -20651
rect 7656 -20703 8019 -20651
rect 8073 -20703 8083 -20650
rect 7656 -20704 8083 -20703
rect 7591 -20715 8083 -20704
rect 12437 -20650 12929 -20639
rect 12437 -20651 12865 -20650
rect 12437 -20704 12448 -20651
rect 12502 -20703 12865 -20651
rect 12919 -20703 12929 -20650
rect 12502 -20704 12929 -20703
rect 12437 -20715 12929 -20704
rect 17283 -20650 17775 -20639
rect 17283 -20651 17711 -20650
rect 17283 -20704 17294 -20651
rect 17348 -20703 17711 -20651
rect 17765 -20703 17775 -20650
rect 17348 -20704 17775 -20703
rect 17283 -20715 17775 -20704
rect 22129 -20650 22621 -20639
rect 22129 -20651 22557 -20650
rect 22129 -20704 22140 -20651
rect 22194 -20703 22557 -20651
rect 22611 -20703 22621 -20650
rect 22194 -20704 22621 -20703
rect 22129 -20715 22621 -20704
rect 26975 -20650 27467 -20639
rect 26975 -20651 27403 -20650
rect 26975 -20704 26986 -20651
rect 27040 -20703 27403 -20651
rect 27457 -20703 27467 -20650
rect 27040 -20704 27467 -20703
rect 26975 -20715 27467 -20704
rect 31821 -20650 32313 -20639
rect 31821 -20651 32249 -20650
rect 31821 -20704 31832 -20651
rect 31886 -20703 32249 -20651
rect 32303 -20703 32313 -20650
rect 31886 -20704 32313 -20703
rect 31821 -20715 32313 -20704
rect 36667 -20650 37159 -20639
rect 36667 -20651 37095 -20650
rect 36667 -20704 36678 -20651
rect 36732 -20703 37095 -20651
rect 37149 -20703 37159 -20650
rect 36732 -20704 37159 -20703
rect 36667 -20715 37159 -20704
rect 7798 -21056 7874 -20715
rect 12644 -21056 12720 -20715
rect 17490 -21056 17566 -20715
rect 22336 -21056 22412 -20715
rect 27182 -21056 27258 -20715
rect 32028 -21056 32104 -20715
rect 36874 -21056 36950 -20715
rect 7392 -21112 42855 -21056
rect 7392 -21168 42672 -21112
rect 42728 -21168 42855 -21112
rect 7392 -21224 42855 -21168
<< via2 >>
rect 3696 2436 3752 2492
rect 8568 2436 8624 2492
rect 13496 2438 13552 2494
rect 18256 2435 18312 2491
rect 23184 2436 23240 2492
rect 28000 2441 28056 2497
rect 32872 2408 32928 2464
rect 37744 2408 37800 2464
rect 13716 1273 13780 1278
rect 13716 1206 13719 1273
rect 13719 1206 13776 1273
rect 13776 1206 13780 1273
rect 13716 1203 13780 1206
rect 18562 1254 18631 1257
rect 18562 1188 18565 1254
rect 18565 1188 18626 1254
rect 18626 1188 18631 1254
rect 18562 1185 18631 1188
rect 23403 1298 23468 1301
rect 23403 1229 23407 1298
rect 23407 1229 23464 1298
rect 23464 1229 23468 1298
rect 23403 1223 23468 1229
rect 28271 1287 28344 1291
rect 28271 1224 28280 1287
rect 28280 1224 28337 1287
rect 28337 1224 28344 1287
rect 28271 1218 28344 1224
rect 33095 1202 33156 1262
rect 6718 883 6790 888
rect 6718 822 6722 883
rect 6722 822 6785 883
rect 6785 822 6790 883
rect 6718 819 6790 822
rect 4029 485 4032 537
rect 4032 485 4088 537
rect 4088 485 4093 537
rect 4029 480 4093 485
rect 3099 -1792 3170 -1736
rect 4033 -15 4092 -13
rect 4033 -67 4035 -15
rect 4035 -67 4089 -15
rect 4089 -67 4092 -15
rect 4033 -69 4092 -67
rect 3696 -983 3700 -907
rect 3700 -983 3768 -907
rect 3768 -983 3774 -907
rect 8880 -14 8938 -12
rect 8880 -66 8882 -14
rect 8882 -66 8934 -14
rect 8934 -66 8938 -14
rect 8880 -68 8938 -66
rect 8574 -983 8632 -907
rect 13725 -15 13784 -13
rect 13725 -67 13727 -15
rect 13727 -67 13782 -15
rect 13782 -67 13784 -15
rect 13725 -69 13784 -67
rect 8391 -1390 8467 -1334
rect 13505 -974 13567 -916
rect 18570 -15 18632 -12
rect 18570 -68 18573 -15
rect 18573 -68 18628 -15
rect 18628 -68 18632 -15
rect 18570 -70 18632 -68
rect 13262 -1389 13338 -1333
rect 18256 -918 18315 -915
rect 18256 -970 18259 -918
rect 18259 -970 18311 -918
rect 18311 -970 18315 -918
rect 18256 -972 18315 -970
rect 18079 -1380 18157 -1324
rect 23418 -14 23476 -12
rect 23418 -67 23420 -14
rect 23420 -67 23474 -14
rect 23474 -67 23476 -14
rect 23418 -69 23476 -67
rect 23194 -916 23260 -913
rect 23194 -968 23199 -916
rect 23199 -968 23256 -916
rect 23256 -968 23260 -916
rect 23194 -971 23260 -968
rect 22962 -1391 23018 -1335
rect 28262 -15 28325 -13
rect 28262 -67 28264 -15
rect 28264 -67 28322 -15
rect 28322 -67 28325 -15
rect 28262 -69 28325 -67
rect 27999 -918 28058 -915
rect 27999 -971 28001 -918
rect 28001 -971 28056 -918
rect 28056 -971 28058 -918
rect 27999 -975 28058 -971
rect 27778 -1390 27834 -1334
rect 33109 -15 33168 -13
rect 33109 -68 33111 -15
rect 33111 -68 33166 -15
rect 33166 -68 33168 -15
rect 33109 -70 33168 -68
rect 32869 -972 32932 -915
rect 32647 -1392 32703 -1336
rect 37744 -971 37800 -915
rect 37492 -1391 37548 -1335
rect 42672 -1568 42728 -1512
rect 3514 -1788 3582 -1722
rect 4895 -1798 4951 -1742
rect 3092 -4607 3148 -4551
rect 4035 -2814 4092 -2812
rect 4035 -2867 4037 -2814
rect 4037 -2867 4090 -2814
rect 4090 -2867 4092 -2814
rect 4035 -2868 4092 -2867
rect 3687 -3783 3755 -3707
rect 9776 -2192 9832 -2136
rect 8879 -2815 8938 -2812
rect 8879 -2867 8882 -2815
rect 8882 -2867 8936 -2815
rect 8936 -2867 8938 -2815
rect 8879 -2870 8938 -2867
rect 8568 -3783 8628 -3707
rect 14584 -2193 14640 -2137
rect 8401 -4187 8457 -4131
rect 13725 -2814 13784 -2812
rect 13725 -2867 13727 -2814
rect 13727 -2867 13782 -2814
rect 13782 -2867 13784 -2814
rect 13725 -2869 13784 -2867
rect 13507 -3717 13570 -3714
rect 13507 -3772 13510 -3717
rect 13510 -3772 13566 -3717
rect 13566 -3772 13570 -3717
rect 13507 -3774 13570 -3772
rect 19463 -2198 19519 -2142
rect 13271 -4188 13327 -4132
rect 18570 -2815 18629 -2812
rect 18570 -2867 18573 -2815
rect 18573 -2867 18627 -2815
rect 18627 -2867 18629 -2815
rect 18570 -2870 18629 -2867
rect 18259 -3719 18323 -3716
rect 18259 -3773 18261 -3719
rect 18261 -3773 18319 -3719
rect 18319 -3773 18323 -3719
rect 18259 -3777 18323 -3773
rect 24273 -2195 24329 -2139
rect 18090 -4178 18146 -4122
rect 23416 -2815 23475 -2813
rect 23416 -2868 23418 -2815
rect 23418 -2868 23472 -2815
rect 23472 -2868 23475 -2815
rect 23416 -2870 23475 -2868
rect 29147 -2196 29203 -2140
rect 23194 -3774 23253 -3718
rect 28265 -2812 28322 -2810
rect 28265 -2866 28267 -2812
rect 28267 -2866 28320 -2812
rect 28320 -2866 28322 -2812
rect 28265 -2868 28322 -2866
rect 22961 -4192 23017 -4136
rect 27990 -3718 28052 -3714
rect 27990 -3770 27993 -3718
rect 27993 -3770 28049 -3718
rect 28049 -3770 28052 -3718
rect 27990 -3772 28052 -3770
rect 33993 -2195 34049 -2139
rect 27777 -4191 27833 -4135
rect 33110 -2815 33166 -2813
rect 33110 -2867 33112 -2815
rect 33112 -2867 33164 -2815
rect 33164 -2867 33166 -2815
rect 33110 -2869 33166 -2867
rect 32869 -3774 32932 -3714
rect 38835 -2195 38891 -2139
rect 32649 -4191 32705 -4135
rect 37744 -3770 37800 -3714
rect 37465 -4192 37521 -4136
rect 42672 -4368 42728 -4312
rect 3472 -4594 3528 -4538
rect 4894 -4595 4950 -4539
rect 3089 -7393 3145 -7337
rect 4035 -5614 4091 -5612
rect 4035 -5666 4037 -5614
rect 4037 -5666 4089 -5614
rect 4089 -5666 4091 -5614
rect 4035 -5668 4091 -5666
rect 3691 -6583 3750 -6507
rect 9775 -4994 9831 -4938
rect 8878 -5615 8937 -5613
rect 8878 -5667 8882 -5615
rect 8882 -5667 8935 -5615
rect 8935 -5667 8937 -5615
rect 8878 -5670 8937 -5667
rect 8565 -6583 8624 -6507
rect 14584 -4997 14640 -4941
rect 8399 -6990 8455 -6934
rect 13725 -5615 13783 -5613
rect 13725 -5667 13728 -5615
rect 13728 -5667 13780 -5615
rect 13780 -5667 13783 -5615
rect 13725 -5669 13783 -5667
rect 13506 -6515 13569 -6513
rect 13506 -6571 13508 -6515
rect 13508 -6571 13566 -6515
rect 13566 -6571 13569 -6515
rect 13506 -6573 13569 -6571
rect 19462 -4993 19518 -4937
rect 13250 -6982 13306 -6926
rect 18569 -5612 18634 -5607
rect 18569 -5667 18574 -5612
rect 18574 -5667 18629 -5612
rect 18629 -5667 18634 -5612
rect 18569 -5671 18634 -5667
rect 18253 -6520 18318 -6517
rect 18253 -6573 18257 -6520
rect 18257 -6573 18315 -6520
rect 18315 -6573 18318 -6520
rect 18253 -6577 18318 -6573
rect 24273 -4990 24329 -4934
rect 18089 -6992 18145 -6936
rect 23416 -5614 23478 -5610
rect 23416 -5667 23420 -5614
rect 23420 -5667 23473 -5614
rect 23473 -5667 23478 -5614
rect 23416 -5671 23478 -5667
rect 23194 -6517 23252 -6516
rect 23194 -6572 23250 -6517
rect 23250 -6572 23252 -6517
rect 29147 -4991 29203 -4935
rect 22960 -6993 23016 -6937
rect 28264 -5614 28323 -5611
rect 28264 -5666 28267 -5614
rect 28267 -5666 28319 -5614
rect 28319 -5666 28323 -5614
rect 28264 -5668 28323 -5666
rect 27985 -6519 28045 -6515
rect 27985 -6574 27989 -6519
rect 27989 -6574 28042 -6519
rect 28042 -6574 28045 -6519
rect 27985 -6576 28045 -6574
rect 33992 -4990 34048 -4934
rect 27773 -6988 27829 -6932
rect 33109 -5614 33169 -5611
rect 33109 -5667 33111 -5614
rect 33111 -5667 33165 -5614
rect 33165 -5667 33169 -5614
rect 33109 -5669 33169 -5667
rect 38833 -5506 38894 -5502
rect 38833 -5558 38894 -5506
rect 32870 -6518 32933 -6517
rect 32870 -6573 32933 -6518
rect 32649 -6990 32705 -6934
rect 37744 -6570 37800 -6514
rect 42671 -7168 42728 -7112
rect 3470 -7393 3526 -7337
rect 4898 -7398 4954 -7342
rect 3302 -10199 3358 -10143
rect 4034 -8415 4091 -8413
rect 4034 -8467 4036 -8415
rect 4036 -8467 4089 -8415
rect 4089 -8467 4091 -8415
rect 4034 -8469 4091 -8467
rect 9775 -7792 9831 -7736
rect 3696 -9373 3752 -9317
rect 8878 -8414 8942 -8411
rect 8878 -8469 8882 -8414
rect 8882 -8469 8938 -8414
rect 8938 -8469 8942 -8414
rect 8878 -8471 8942 -8469
rect 8566 -9383 8627 -9307
rect 14584 -7789 14640 -7733
rect 8401 -9791 8457 -9735
rect 13726 -8415 13782 -8413
rect 13726 -8467 13728 -8415
rect 13728 -8467 13780 -8415
rect 13780 -8467 13782 -8415
rect 13726 -8469 13782 -8467
rect 13505 -9316 13570 -9314
rect 13505 -9371 13510 -9316
rect 13510 -9371 13567 -9316
rect 13567 -9371 13570 -9316
rect 13505 -9373 13570 -9371
rect 19462 -7792 19518 -7736
rect 13245 -9788 13301 -9732
rect 18571 -8470 18629 -8412
rect 18252 -9321 18318 -9317
rect 18252 -9373 18256 -9321
rect 18256 -9373 18314 -9321
rect 18314 -9373 18318 -9321
rect 18252 -9376 18318 -9373
rect 24273 -7793 24329 -7737
rect 18088 -9790 18144 -9734
rect 23416 -8413 23479 -8406
rect 23416 -8468 23420 -8413
rect 23420 -8468 23475 -8413
rect 23475 -8468 23479 -8413
rect 23416 -8471 23479 -8468
rect 23194 -9316 23252 -9314
rect 23194 -9371 23196 -9316
rect 23196 -9371 23250 -9316
rect 23250 -9371 23252 -9316
rect 23194 -9373 23252 -9371
rect 29149 -7790 29205 -7734
rect 22961 -9796 23017 -9740
rect 28262 -8413 28323 -8411
rect 28262 -8467 28264 -8413
rect 28264 -8467 28321 -8413
rect 28321 -8467 28323 -8413
rect 28262 -8469 28323 -8467
rect 27993 -9375 28053 -9317
rect 33993 -7790 34049 -7734
rect 27778 -9793 27834 -9737
rect 33107 -8414 33166 -8413
rect 33107 -8469 33110 -8414
rect 33110 -8469 33165 -8414
rect 33165 -8469 33166 -8414
rect 33107 -8471 33166 -8469
rect 38833 -7794 38889 -7738
rect 32867 -9317 32933 -9316
rect 32867 -9372 32868 -9317
rect 32868 -9372 32932 -9317
rect 32932 -9372 32933 -9317
rect 32867 -9374 32933 -9372
rect 32646 -9795 32702 -9739
rect 37744 -9371 37800 -9315
rect 37465 -9792 37521 -9736
rect 42672 -9968 42728 -9912
rect 3473 -10194 3529 -10138
rect 4896 -10200 4952 -10144
rect 4035 -11214 4091 -11212
rect 4035 -11266 4037 -11214
rect 4037 -11266 4089 -11214
rect 4089 -11266 4091 -11214
rect 4035 -11268 4091 -11266
rect 3205 -13001 3261 -12945
rect 3688 -12183 3758 -12107
rect 9776 -10590 9832 -10534
rect 8874 -11272 8938 -11212
rect 8559 -12118 8617 -12114
rect 8559 -12171 8562 -12118
rect 8562 -12171 8614 -12118
rect 8614 -12171 8617 -12118
rect 8559 -12174 8617 -12171
rect 14584 -10591 14640 -10535
rect 8401 -12589 8457 -12533
rect 13726 -11214 13782 -11212
rect 13726 -11266 13728 -11214
rect 13728 -11266 13780 -11214
rect 13780 -11266 13782 -11214
rect 13726 -11269 13782 -11266
rect 13504 -12119 13564 -12116
rect 13504 -12171 13506 -12119
rect 13506 -12171 13560 -12119
rect 13560 -12171 13564 -12119
rect 13504 -12173 13564 -12171
rect 19462 -10591 19518 -10535
rect 13250 -12585 13306 -12529
rect 18571 -11213 18630 -11210
rect 18571 -11268 18573 -11213
rect 18573 -11268 18626 -11213
rect 18626 -11268 18630 -11213
rect 18571 -11270 18630 -11268
rect 18249 -12121 18313 -12118
rect 18249 -12174 18253 -12121
rect 18253 -12174 18309 -12121
rect 18309 -12174 18313 -12121
rect 18249 -12177 18313 -12174
rect 24274 -10590 24330 -10534
rect 18092 -12589 18148 -12533
rect 23417 -11213 23480 -11210
rect 23417 -11267 23420 -11213
rect 23420 -11267 23477 -11213
rect 23477 -11267 23480 -11213
rect 23417 -11270 23480 -11267
rect 23190 -12116 23255 -12113
rect 23190 -12173 23192 -12116
rect 23192 -12173 23252 -12116
rect 23252 -12173 23255 -12116
rect 23190 -12176 23255 -12173
rect 29147 -10589 29203 -10533
rect 22932 -12593 22988 -12537
rect 28264 -11214 28320 -11212
rect 28264 -11266 28266 -11214
rect 28266 -11266 28318 -11214
rect 28318 -11266 28320 -11214
rect 28264 -11268 28320 -11266
rect 33992 -10592 34048 -10536
rect 27998 -12175 28058 -12117
rect 27776 -12589 27832 -12533
rect 33111 -11216 33167 -11212
rect 33111 -11268 33164 -11216
rect 33164 -11268 33167 -11216
rect 38836 -10590 38892 -10534
rect 32888 -12119 32944 -12116
rect 32888 -12171 32889 -12119
rect 32889 -12171 32941 -12119
rect 32941 -12171 32944 -12119
rect 32888 -12173 32944 -12171
rect 32648 -12592 32704 -12536
rect 37744 -12170 37800 -12114
rect 37466 -12590 37522 -12534
rect 42672 -12768 42728 -12712
rect 3469 -12996 3525 -12940
rect 4895 -12996 4951 -12940
rect 4035 -14015 4092 -14013
rect 4035 -14067 4037 -14015
rect 4037 -14067 4089 -14015
rect 4089 -14067 4092 -14015
rect 4035 -14070 4092 -14067
rect 3191 -15794 3247 -15738
rect 3681 -14983 3746 -14907
rect 9774 -13396 9830 -13340
rect 8879 -14013 8939 -14011
rect 8879 -14067 8882 -14013
rect 8882 -14067 8937 -14013
rect 8937 -14067 8939 -14013
rect 8879 -14069 8939 -14067
rect 8578 -14919 8636 -14917
rect 8578 -14971 8581 -14919
rect 8581 -14971 8633 -14919
rect 8633 -14971 8636 -14919
rect 8578 -14973 8636 -14971
rect 14583 -13391 14639 -13335
rect 8402 -15393 8458 -15337
rect 13725 -14014 13784 -14012
rect 13725 -14067 13727 -14014
rect 13727 -14067 13782 -14014
rect 13782 -14067 13784 -14014
rect 13725 -14069 13784 -14067
rect 13509 -14918 13568 -14916
rect 13509 -14971 13512 -14918
rect 13512 -14971 13567 -14918
rect 13567 -14971 13568 -14918
rect 13509 -14973 13568 -14971
rect 19461 -13389 19517 -13333
rect 13248 -15395 13304 -15339
rect 18572 -14013 18630 -14011
rect 18572 -14068 18630 -14013
rect 18252 -14921 18316 -14917
rect 18252 -14974 18256 -14921
rect 18256 -14974 18312 -14921
rect 18312 -14974 18316 -14921
rect 18252 -14979 18316 -14974
rect 24275 -13390 24331 -13334
rect 18091 -15391 18147 -15335
rect 23417 -14015 23477 -14013
rect 23417 -14068 23419 -14015
rect 23419 -14068 23474 -14015
rect 23474 -14068 23477 -14015
rect 23417 -14070 23477 -14068
rect 23191 -14913 23254 -14909
rect 23191 -14971 23196 -14913
rect 23196 -14971 23251 -14913
rect 23251 -14971 23254 -14913
rect 23191 -14974 23254 -14971
rect 29148 -13388 29204 -13332
rect 22960 -15391 23016 -15335
rect 28263 -14013 28321 -14012
rect 28263 -14067 28264 -14013
rect 28264 -14067 28320 -14013
rect 28320 -14067 28321 -14013
rect 28263 -14068 28321 -14067
rect 33993 -13391 34049 -13335
rect 27997 -14972 28062 -14916
rect 27777 -15391 27833 -15335
rect 33110 -14014 33166 -14012
rect 33110 -14067 33112 -14014
rect 33112 -14067 33164 -14014
rect 33164 -14067 33166 -14014
rect 33110 -14069 33166 -14067
rect 38837 -13391 38893 -13335
rect 32866 -14918 32938 -14916
rect 32866 -14973 32868 -14918
rect 32868 -14973 32936 -14918
rect 32936 -14973 32938 -14918
rect 32866 -14974 32938 -14973
rect 32648 -15388 32704 -15332
rect 37744 -14970 37800 -14914
rect 37464 -15387 37520 -15331
rect 42672 -15568 42728 -15512
rect 3471 -15802 3527 -15746
rect 4898 -15796 4954 -15740
rect 4034 -16815 4090 -16812
rect 4034 -16867 4036 -16815
rect 4036 -16867 4088 -16815
rect 4088 -16867 4090 -16815
rect 4034 -16868 4090 -16867
rect 3692 -17783 3760 -17707
rect 9774 -16196 9830 -16140
rect 8879 -16815 8938 -16812
rect 8879 -16867 8882 -16815
rect 8882 -16867 8934 -16815
rect 8934 -16867 8938 -16815
rect 8879 -16870 8938 -16867
rect 8570 -17720 8630 -17717
rect 8570 -17772 8572 -17720
rect 8572 -17772 8626 -17720
rect 8626 -17772 8630 -17720
rect 8570 -17775 8630 -17772
rect 14584 -16193 14640 -16137
rect 8400 -18193 8456 -18137
rect 13726 -16814 13785 -16812
rect 13726 -16867 13728 -16814
rect 13728 -16867 13783 -16814
rect 13783 -16867 13785 -16814
rect 13726 -16869 13785 -16867
rect 19463 -16191 19519 -16135
rect 13505 -17717 13561 -17715
rect 13505 -17769 13507 -17717
rect 13507 -17769 13559 -17717
rect 13559 -17769 13561 -17717
rect 13505 -17771 13561 -17769
rect 13262 -18196 13318 -18140
rect 18572 -16814 18630 -16810
rect 18572 -16868 18573 -16814
rect 18573 -16868 18627 -16814
rect 18627 -16868 18630 -16814
rect 18572 -16869 18630 -16868
rect 18250 -17717 18318 -17715
rect 18250 -17773 18253 -17717
rect 18253 -17773 18315 -17717
rect 18315 -17773 18318 -17717
rect 18250 -17776 18318 -17773
rect 24273 -16198 24329 -16142
rect 18090 -18190 18146 -18134
rect 23415 -16814 23478 -16811
rect 23415 -16867 23419 -16814
rect 23419 -16867 23475 -16814
rect 23475 -16867 23478 -16814
rect 23415 -16870 23478 -16867
rect 23191 -17714 23251 -17712
rect 23191 -17775 23197 -17714
rect 23197 -17775 23250 -17714
rect 23250 -17775 23251 -17714
rect 23191 -17778 23251 -17775
rect 29148 -16190 29204 -16134
rect 22956 -18190 23012 -18134
rect 28265 -16814 28323 -16811
rect 28265 -16866 28267 -16814
rect 28267 -16866 28320 -16814
rect 28320 -16866 28323 -16814
rect 28265 -16867 28323 -16866
rect 27999 -17716 28060 -17712
rect 27999 -17769 28060 -17716
rect 33993 -16190 34049 -16134
rect 27779 -18192 27835 -18136
rect 33109 -16815 33167 -16813
rect 33109 -16867 33112 -16815
rect 33112 -16867 33165 -16815
rect 33165 -16867 33167 -16815
rect 33109 -16870 33167 -16867
rect 38835 -16191 38891 -16135
rect 32868 -17775 32935 -17715
rect 32646 -18194 32702 -18138
rect 37744 -17772 37800 -17716
rect 42672 -18368 42728 -18312
rect 3471 -18569 3527 -18513
rect 4893 -19502 4956 -19499
rect 4893 -19555 4956 -19502
rect 4034 -19615 4091 -19613
rect 4034 -19668 4036 -19615
rect 4036 -19668 4089 -19615
rect 4089 -19668 4091 -19615
rect 4034 -19669 4091 -19668
rect 3696 -20583 3752 -20507
rect 9772 -19501 9834 -19498
rect 9772 -19554 9834 -19501
rect 8881 -19614 8939 -19612
rect 8881 -19666 8882 -19614
rect 8882 -19666 8936 -19614
rect 8936 -19666 8939 -19614
rect 8881 -19668 8939 -19666
rect 8563 -20518 8625 -20514
rect 8563 -20570 8568 -20518
rect 8568 -20570 8620 -20518
rect 8620 -20570 8625 -20518
rect 8563 -20573 8625 -20570
rect 14580 -19505 14645 -19501
rect 14580 -19557 14645 -19505
rect 13727 -19614 13784 -19612
rect 13727 -19666 13729 -19614
rect 13729 -19666 13781 -19614
rect 13781 -19666 13784 -19614
rect 13727 -19668 13784 -19666
rect 19458 -19506 19521 -19502
rect 19458 -19558 19521 -19506
rect 18573 -19669 18630 -19613
rect 13513 -20518 13571 -20515
rect 13513 -20570 13515 -20518
rect 13515 -20570 13568 -20518
rect 13568 -20570 13571 -20518
rect 13513 -20571 13571 -20570
rect 18251 -20521 18315 -20518
rect 18251 -20577 18254 -20521
rect 18254 -20577 18312 -20521
rect 18312 -20577 18315 -20521
rect 18251 -20580 18315 -20577
rect 24269 -19503 24334 -19499
rect 24269 -19556 24334 -19503
rect 23417 -19615 23476 -19612
rect 23417 -19667 23419 -19615
rect 23419 -19667 23474 -19615
rect 23474 -19667 23476 -19615
rect 23417 -19669 23476 -19667
rect 23193 -20517 23253 -20514
rect 23193 -20574 23198 -20517
rect 23198 -20574 23250 -20517
rect 23250 -20574 23253 -20517
rect 23193 -20577 23253 -20574
rect 29145 -19505 29206 -19502
rect 29145 -19558 29206 -19505
rect 28262 -19614 28319 -19612
rect 28262 -19667 28263 -19614
rect 28263 -19667 28318 -19614
rect 28318 -19667 28319 -19614
rect 28262 -19669 28319 -19667
rect 27998 -20574 28059 -20517
rect 33989 -19505 34051 -19501
rect 33989 -19557 34051 -19505
rect 33108 -19614 33170 -19611
rect 33108 -19668 33111 -19614
rect 33111 -19668 33166 -19614
rect 33166 -19668 33170 -19614
rect 33108 -19670 33170 -19668
rect 32869 -20574 32932 -20517
rect 42672 -21168 42728 -21112
<< metal3 >>
rect 3686 2492 3762 2502
rect 3686 2436 3696 2492
rect 3752 2436 3762 2492
rect 3686 2426 3762 2436
rect 8558 2492 8634 2502
rect 8558 2436 8568 2492
rect 8624 2436 8634 2492
rect 8558 2426 8634 2436
rect 13486 2494 13562 2504
rect 13486 2438 13496 2494
rect 13552 2438 13562 2494
rect 13486 2428 13562 2438
rect 18246 2491 18322 2501
rect 18246 2435 18256 2491
rect 18312 2435 18322 2491
rect 18246 2425 18322 2435
rect 23174 2492 23250 2502
rect 23174 2436 23184 2492
rect 23240 2436 23250 2492
rect 23174 2426 23250 2436
rect 27987 2497 28069 2509
rect 27987 2441 28000 2497
rect 28056 2441 28069 2497
rect 27987 2429 28069 2441
rect 32858 2464 32939 2476
rect 32858 2408 32872 2464
rect 32928 2408 32939 2464
rect 32858 2394 32939 2408
rect 37734 2464 37810 2474
rect 37734 2408 37744 2464
rect 37800 2408 37810 2464
rect 37734 2398 37810 2408
rect 23370 1301 23497 1314
rect 13688 1278 13804 1299
rect 13688 1203 13716 1278
rect 13780 1203 13804 1278
rect 13688 1181 13804 1203
rect 18536 1257 18648 1264
rect 18536 1185 18562 1257
rect 18631 1185 18648 1257
rect 23370 1223 23403 1301
rect 23468 1223 23497 1301
rect 23370 1196 23497 1223
rect 28247 1291 28370 1304
rect 28247 1218 28271 1291
rect 28344 1218 28370 1291
rect 28247 1192 28370 1218
rect 33065 1262 33188 1274
rect 33065 1202 33095 1262
rect 33156 1202 33188 1262
rect 18536 1166 18648 1185
rect 33065 1176 33188 1202
rect 6693 888 6807 894
rect 6693 819 6718 888
rect 6790 880 6807 888
rect 6790 876 8945 880
rect 6790 819 8856 876
rect 6693 813 8856 819
rect 8928 813 8945 876
rect 6693 808 8945 813
rect 6693 804 6807 808
rect 3998 537 4115 539
rect 3998 480 4029 537
rect 4093 480 4115 537
rect 3998 448 4115 480
rect 4010 -13 4115 -1
rect 4010 -69 4033 -13
rect 4092 -69 4115 -13
rect 4010 -78 4115 -69
rect 8859 -12 8951 -8
rect 8859 -68 8880 -12
rect 8938 -68 8951 -12
rect 8859 -74 8951 -68
rect 13701 -13 13810 -1
rect 13701 -69 13725 -13
rect 13784 -69 13810 -13
rect 13701 -78 13810 -69
rect 18553 -12 18646 2
rect 18553 -70 18570 -12
rect 18632 -70 18646 -12
rect 18553 -84 18646 -70
rect 23405 -12 23487 -1
rect 23405 -69 23418 -12
rect 23476 -69 23487 -12
rect 23405 -80 23487 -69
rect 28249 -13 28338 1
rect 28249 -69 28262 -13
rect 28325 -69 28338 -13
rect 28249 -83 28338 -69
rect 33097 -13 33182 -3
rect 33097 -70 33109 -13
rect 33168 -70 33182 -13
rect 33097 -79 33182 -70
rect 3672 -907 3794 -884
rect 3672 -983 3696 -907
rect 3774 -983 3794 -907
rect 3672 -1002 3794 -983
rect 8545 -907 8658 -893
rect 8545 -983 8574 -907
rect 8632 -983 8658 -907
rect 8545 -1000 8658 -983
rect 13469 -916 13581 -896
rect 13469 -974 13505 -916
rect 13567 -974 13581 -916
rect 13469 -998 13581 -974
rect 18223 -915 18325 -896
rect 18223 -972 18256 -915
rect 18315 -972 18325 -915
rect 18223 -996 18325 -972
rect 23156 -913 23270 -895
rect 23156 -971 23194 -913
rect 23260 -971 23270 -913
rect 23156 -999 23270 -971
rect 27975 -915 28081 -898
rect 27975 -975 27999 -915
rect 28058 -975 28081 -915
rect 27975 -1001 28081 -975
rect 32850 -915 32947 -897
rect 32850 -972 32869 -915
rect 32932 -972 32947 -915
rect 32850 -990 32947 -972
rect 37732 -915 37811 -905
rect 37732 -971 37744 -915
rect 37800 -971 37811 -915
rect 37732 -981 37811 -971
rect 8391 -1334 8467 -1324
rect 3460 -1680 3536 -1679
rect 8391 -1680 8467 -1390
rect 13262 -1333 13338 -1323
rect 13262 -1680 13338 -1389
rect 18079 -1324 18157 -1314
rect 18079 -1402 18157 -1380
rect 22952 -1335 23028 -1325
rect 22952 -1391 22962 -1335
rect 23018 -1391 23028 -1335
rect 18079 -1680 18155 -1402
rect 22952 -1680 23028 -1391
rect 27766 -1334 27842 -1324
rect 27766 -1390 27778 -1334
rect 27834 -1390 27842 -1334
rect 37482 -1335 37558 -1325
rect 27766 -1680 27842 -1390
rect 32637 -1392 32647 -1336
rect 32703 -1392 32713 -1336
rect 32637 -1680 32713 -1392
rect 37482 -1391 37492 -1335
rect 37548 -1391 37558 -1335
rect 37482 -1680 37558 -1391
rect 42662 -1512 42738 -1502
rect 42662 -1568 42672 -1512
rect 42728 -1568 42738 -1512
rect 42662 -1578 42738 -1568
rect 3024 -1722 39032 -1680
rect 3024 -1736 3514 -1722
rect 3024 -1792 3099 -1736
rect 3170 -1788 3514 -1736
rect 3582 -1742 39032 -1722
rect 3582 -1788 4895 -1742
rect 3170 -1792 4895 -1788
rect 3024 -1798 4895 -1792
rect 4951 -1798 39032 -1742
rect 3024 -1848 39032 -1798
rect 9762 -2136 9844 -1848
rect 9762 -2192 9776 -2136
rect 9832 -2192 9844 -2136
rect 14570 -2137 14655 -1848
rect 14570 -2193 14584 -2137
rect 14640 -2193 14655 -2137
rect 19448 -2142 19531 -1848
rect 19448 -2198 19463 -2142
rect 19519 -2198 19531 -2142
rect 24259 -2139 24344 -1848
rect 24259 -2195 24273 -2139
rect 24329 -2195 24344 -2139
rect 24259 -2205 24344 -2195
rect 29135 -2140 29216 -1848
rect 29135 -2196 29147 -2140
rect 29203 -2196 29216 -2140
rect 33979 -2139 34061 -1848
rect 33979 -2195 33993 -2139
rect 34049 -2195 34061 -2139
rect 38823 -2139 38903 -1848
rect 38823 -2195 38835 -2139
rect 38891 -2195 38903 -2139
rect 29135 -2206 29216 -2196
rect 38823 -2205 38903 -2195
rect 4009 -2812 4115 -2806
rect 4009 -2868 4035 -2812
rect 4092 -2868 4115 -2812
rect 4009 -2875 4115 -2868
rect 8860 -2812 8959 -2807
rect 8860 -2870 8879 -2812
rect 8938 -2870 8959 -2812
rect 8860 -2876 8959 -2870
rect 13704 -2812 13805 -2804
rect 13704 -2869 13725 -2812
rect 13784 -2869 13805 -2812
rect 13704 -2882 13805 -2869
rect 18558 -2812 18642 -2798
rect 18558 -2870 18570 -2812
rect 18629 -2870 18642 -2812
rect 18558 -2878 18642 -2870
rect 23402 -2813 23491 -2796
rect 23402 -2870 23416 -2813
rect 23475 -2870 23491 -2813
rect 23402 -2883 23491 -2870
rect 28246 -2810 28340 -2801
rect 28246 -2868 28265 -2810
rect 28322 -2868 28340 -2810
rect 28246 -2881 28340 -2868
rect 33092 -2813 33180 -2801
rect 33092 -2869 33110 -2813
rect 33166 -2869 33180 -2813
rect 33092 -2880 33180 -2869
rect 3655 -3707 3779 -3692
rect 3655 -3783 3687 -3707
rect 3755 -3783 3779 -3707
rect 3655 -3800 3779 -3783
rect 8539 -3707 8643 -3693
rect 8539 -3783 8568 -3707
rect 8628 -3783 8643 -3707
rect 8539 -3797 8643 -3783
rect 13472 -3714 13586 -3692
rect 13472 -3774 13507 -3714
rect 13570 -3774 13586 -3714
rect 13472 -3803 13586 -3774
rect 18233 -3716 18335 -3695
rect 18233 -3777 18259 -3716
rect 18323 -3777 18335 -3716
rect 18233 -3801 18335 -3777
rect 23155 -3718 23270 -3699
rect 23155 -3774 23194 -3718
rect 23253 -3774 23270 -3718
rect 23155 -3796 23270 -3774
rect 27965 -3714 28068 -3696
rect 27965 -3772 27990 -3714
rect 28052 -3772 28068 -3714
rect 27965 -3796 28068 -3772
rect 32843 -3714 32940 -3695
rect 32843 -3774 32869 -3714
rect 32932 -3774 32940 -3714
rect 32843 -3788 32940 -3774
rect 37731 -3714 37810 -3704
rect 37731 -3770 37744 -3714
rect 37800 -3770 37810 -3714
rect 37731 -3780 37810 -3770
rect 8391 -4131 8467 -4130
rect 8391 -4187 8401 -4131
rect 8457 -4187 8467 -4131
rect 3054 -4480 3190 -4479
rect 8391 -4480 8467 -4187
rect 13261 -4188 13271 -4132
rect 13327 -4188 13337 -4132
rect 13261 -4480 13337 -4188
rect 18080 -4178 18090 -4122
rect 18146 -4178 18156 -4122
rect 18080 -4480 18156 -4178
rect 22951 -4136 23027 -4126
rect 22951 -4192 22961 -4136
rect 23017 -4192 23027 -4136
rect 22951 -4480 23027 -4192
rect 27767 -4191 27777 -4135
rect 27833 -4191 27843 -4135
rect 27767 -4480 27843 -4191
rect 32639 -4191 32649 -4135
rect 32705 -4191 32715 -4135
rect 32639 -4480 32715 -4191
rect 37455 -4192 37465 -4136
rect 37521 -4192 37531 -4136
rect 37455 -4480 37531 -4192
rect 42662 -4312 42738 -4302
rect 42662 -4368 42672 -4312
rect 42728 -4368 42738 -4312
rect 42662 -4378 42738 -4368
rect 3024 -4538 39032 -4480
rect 3024 -4551 3472 -4538
rect 3024 -4607 3092 -4551
rect 3148 -4594 3472 -4551
rect 3528 -4539 39032 -4538
rect 3528 -4594 4894 -4539
rect 3148 -4595 4894 -4594
rect 4950 -4595 39032 -4539
rect 3148 -4607 39032 -4595
rect 3024 -4648 39032 -4607
rect 3054 -4649 3190 -4648
rect 9762 -4938 9844 -4648
rect 9762 -4994 9775 -4938
rect 9831 -4994 9844 -4938
rect 14570 -4941 14655 -4648
rect 14570 -4997 14584 -4941
rect 14640 -4997 14655 -4941
rect 19448 -4937 19531 -4648
rect 19448 -4993 19462 -4937
rect 19518 -4993 19531 -4937
rect 24259 -4934 24344 -4648
rect 24259 -4990 24273 -4934
rect 24329 -4990 24344 -4934
rect 29135 -4935 29216 -4648
rect 29135 -4991 29147 -4935
rect 29203 -4991 29216 -4935
rect 33979 -4934 34061 -4648
rect 33979 -4990 33992 -4934
rect 34048 -4990 34061 -4934
rect 38823 -5502 38903 -4648
rect 38823 -5558 38833 -5502
rect 38894 -5558 38904 -5502
rect 38823 -5561 38904 -5558
rect 4015 -5612 4108 -5609
rect 4015 -5668 4035 -5612
rect 4091 -5668 4108 -5612
rect 4015 -5675 4108 -5668
rect 8860 -5613 8955 -5608
rect 8860 -5670 8878 -5613
rect 8937 -5670 8955 -5613
rect 8860 -5674 8955 -5670
rect 13701 -5613 13802 -5602
rect 13701 -5669 13725 -5613
rect 13783 -5669 13802 -5613
rect 13701 -5679 13802 -5669
rect 18556 -5607 18645 -5598
rect 18556 -5671 18569 -5607
rect 18634 -5671 18645 -5607
rect 18556 -5682 18645 -5671
rect 23404 -5610 23490 -5601
rect 23404 -5671 23416 -5610
rect 23478 -5671 23490 -5610
rect 23404 -5683 23490 -5671
rect 28251 -5611 28335 -5601
rect 28251 -5668 28264 -5611
rect 28323 -5668 28335 -5611
rect 28251 -5683 28335 -5668
rect 33096 -5611 33179 -5606
rect 33096 -5669 33109 -5611
rect 33169 -5669 33179 -5611
rect 33096 -5679 33179 -5669
rect 3660 -6507 3762 -6493
rect 3660 -6583 3691 -6507
rect 3750 -6583 3762 -6507
rect 3660 -6600 3762 -6583
rect 8529 -6507 8634 -6496
rect 8529 -6583 8565 -6507
rect 8624 -6583 8634 -6507
rect 8529 -6597 8634 -6583
rect 13470 -6513 13579 -6495
rect 13470 -6573 13506 -6513
rect 13569 -6573 13579 -6513
rect 13470 -6597 13579 -6573
rect 18230 -6517 18333 -6492
rect 18230 -6577 18253 -6517
rect 18318 -6577 18333 -6517
rect 18230 -6599 18333 -6577
rect 23153 -6516 23268 -6495
rect 23153 -6572 23194 -6516
rect 23252 -6572 23268 -6516
rect 23153 -6597 23268 -6572
rect 27963 -6515 28073 -6494
rect 27963 -6576 27985 -6515
rect 28045 -6576 28073 -6515
rect 27963 -6597 28073 -6576
rect 32851 -6517 32944 -6500
rect 32851 -6573 32870 -6517
rect 32933 -6573 32944 -6517
rect 32851 -6588 32944 -6573
rect 37733 -6514 37811 -6503
rect 37733 -6570 37744 -6514
rect 37800 -6570 37811 -6514
rect 37733 -6580 37811 -6570
rect 8389 -6990 8399 -6934
rect 8455 -6990 8465 -6934
rect 8389 -7280 8465 -6990
rect 13240 -6982 13250 -6926
rect 13306 -6982 13316 -6926
rect 13240 -7280 13316 -6982
rect 18079 -6992 18089 -6936
rect 18145 -6992 18155 -6936
rect 18079 -7280 18155 -6992
rect 22950 -6993 22960 -6937
rect 23016 -6993 23026 -6937
rect 22950 -7280 23026 -6993
rect 27763 -6988 27773 -6932
rect 27829 -6988 27839 -6932
rect 27763 -7280 27839 -6988
rect 32639 -6990 32649 -6934
rect 32705 -6990 32715 -6934
rect 32639 -7280 32715 -6990
rect 37454 -7280 37530 -7000
rect 42661 -7112 42739 -7102
rect 42661 -7168 42671 -7112
rect 42728 -7168 42739 -7112
rect 42661 -7178 42739 -7168
rect 3024 -7337 39032 -7280
rect 3024 -7393 3089 -7337
rect 3145 -7393 3470 -7337
rect 3526 -7342 39032 -7337
rect 3526 -7393 4898 -7342
rect 3024 -7398 4898 -7393
rect 4954 -7398 39032 -7342
rect 3024 -7448 39032 -7398
rect 9762 -7498 9845 -7448
rect 9762 -7736 9844 -7498
rect 9762 -7792 9775 -7736
rect 9831 -7792 9844 -7736
rect 14570 -7733 14655 -7448
rect 14570 -7789 14584 -7733
rect 14640 -7789 14655 -7733
rect 19448 -7488 19533 -7448
rect 19448 -7736 19531 -7488
rect 19448 -7792 19462 -7736
rect 19518 -7792 19531 -7736
rect 24259 -7737 24344 -7448
rect 27763 -7449 27839 -7448
rect 24259 -7793 24273 -7737
rect 24329 -7793 24344 -7737
rect 29135 -7483 29220 -7448
rect 33979 -7481 34064 -7448
rect 29135 -7734 29216 -7483
rect 29135 -7790 29149 -7734
rect 29205 -7790 29216 -7734
rect 33979 -7734 34061 -7481
rect 33979 -7790 33993 -7734
rect 34049 -7790 34061 -7734
rect 38823 -7483 38908 -7448
rect 38823 -7738 38903 -7483
rect 38823 -7794 38833 -7738
rect 38889 -7794 38903 -7738
rect 4013 -8413 4113 -8406
rect 4013 -8469 4034 -8413
rect 4091 -8469 4113 -8413
rect 4013 -8478 4113 -8469
rect 8854 -8411 8968 -8405
rect 8854 -8471 8878 -8411
rect 8942 -8471 8968 -8411
rect 8854 -8481 8968 -8471
rect 13705 -8413 13804 -8401
rect 13705 -8469 13726 -8413
rect 13782 -8469 13804 -8413
rect 13705 -8478 13804 -8469
rect 18550 -8412 18647 -8398
rect 18550 -8470 18571 -8412
rect 18629 -8470 18647 -8412
rect 18550 -8493 18647 -8470
rect 23405 -8406 23490 -8393
rect 23405 -8471 23416 -8406
rect 23479 -8471 23490 -8406
rect 23405 -8481 23490 -8471
rect 28247 -8411 28343 -8401
rect 28247 -8469 28262 -8411
rect 28323 -8469 28343 -8411
rect 28247 -8487 28343 -8469
rect 33093 -8413 33183 -8403
rect 33093 -8471 33107 -8413
rect 33166 -8471 33183 -8413
rect 33093 -8484 33183 -8471
rect 3670 -9317 3776 -9299
rect 3670 -9373 3696 -9317
rect 3752 -9373 3776 -9317
rect 3670 -9397 3776 -9373
rect 8529 -9307 8645 -9296
rect 8529 -9383 8566 -9307
rect 8627 -9383 8645 -9307
rect 8529 -9402 8645 -9383
rect 13467 -9314 13579 -9296
rect 13467 -9373 13505 -9314
rect 13570 -9373 13579 -9314
rect 13467 -9399 13579 -9373
rect 18226 -9317 18333 -9296
rect 18226 -9376 18252 -9317
rect 18318 -9376 18333 -9317
rect 18226 -9396 18333 -9376
rect 23153 -9314 23265 -9295
rect 23153 -9373 23194 -9314
rect 23252 -9373 23265 -9314
rect 23153 -9397 23265 -9373
rect 27968 -9317 28077 -9293
rect 27968 -9375 27993 -9317
rect 28053 -9375 28077 -9317
rect 27968 -9397 28077 -9375
rect 32853 -9316 32946 -9300
rect 32853 -9374 32867 -9316
rect 32933 -9374 32946 -9316
rect 32853 -9387 32946 -9374
rect 37734 -9315 37811 -9303
rect 37734 -9371 37744 -9315
rect 37800 -9371 37811 -9315
rect 37734 -9381 37811 -9371
rect 13236 -9732 13313 -9725
rect 8391 -9791 8401 -9735
rect 8457 -9791 8467 -9735
rect 8391 -10080 8467 -9791
rect 13236 -9788 13245 -9732
rect 13301 -9788 13313 -9732
rect 13236 -9797 13313 -9788
rect 18078 -9790 18088 -9734
rect 18144 -9790 18154 -9734
rect 13236 -10080 13312 -9797
rect 18078 -10080 18154 -9790
rect 22951 -9796 22961 -9740
rect 23017 -9796 23027 -9740
rect 22951 -10080 23027 -9796
rect 27768 -9793 27778 -9737
rect 27834 -9793 27844 -9737
rect 27768 -10080 27844 -9793
rect 32636 -9795 32646 -9739
rect 32702 -9795 32712 -9739
rect 32636 -10080 32712 -9795
rect 37455 -9792 37465 -9736
rect 37521 -9792 37531 -9736
rect 37455 -10080 37531 -9792
rect 42662 -9912 42738 -9902
rect 42662 -9968 42672 -9912
rect 42728 -9968 42738 -9912
rect 42662 -9978 42738 -9968
rect 3192 -10138 39032 -10080
rect 3192 -10143 3473 -10138
rect 3192 -10199 3302 -10143
rect 3358 -10194 3473 -10143
rect 3529 -10144 39032 -10138
rect 3529 -10194 4896 -10144
rect 3358 -10199 4896 -10194
rect 3192 -10200 4896 -10199
rect 4952 -10200 39032 -10144
rect 3192 -10248 39032 -10200
rect 9762 -10298 9845 -10248
rect 9762 -10534 9844 -10298
rect 9762 -10590 9776 -10534
rect 9832 -10590 9844 -10534
rect 14570 -10535 14655 -10248
rect 14570 -10591 14584 -10535
rect 14640 -10591 14655 -10535
rect 19448 -10288 19533 -10248
rect 19448 -10535 19531 -10288
rect 19448 -10591 19462 -10535
rect 19518 -10591 19531 -10535
rect 24259 -10534 24344 -10248
rect 24259 -10590 24274 -10534
rect 24330 -10590 24344 -10534
rect 29135 -10283 29220 -10248
rect 33979 -10281 34064 -10248
rect 29135 -10533 29216 -10283
rect 29135 -10589 29147 -10533
rect 29203 -10589 29216 -10533
rect 33979 -10536 34061 -10281
rect 24259 -10591 24344 -10590
rect 33979 -10592 33992 -10536
rect 34048 -10592 34061 -10536
rect 38823 -10534 38903 -10248
rect 38823 -10590 38836 -10534
rect 38892 -10590 38903 -10534
rect 4013 -11212 4108 -11207
rect 4013 -11268 4035 -11212
rect 4091 -11268 4108 -11212
rect 4013 -11277 4108 -11268
rect 8855 -11212 8956 -11201
rect 8855 -11272 8874 -11212
rect 8938 -11272 8956 -11212
rect 8855 -11284 8956 -11272
rect 13707 -11212 13797 -11202
rect 13707 -11269 13726 -11212
rect 13782 -11269 13797 -11212
rect 13707 -11284 13797 -11269
rect 18556 -11210 18647 -11195
rect 18556 -11270 18571 -11210
rect 18630 -11270 18647 -11210
rect 18556 -11284 18647 -11270
rect 23405 -11210 23490 -11197
rect 23405 -11270 23417 -11210
rect 23480 -11270 23490 -11210
rect 23405 -11283 23490 -11270
rect 28248 -11212 28335 -11204
rect 28248 -11268 28264 -11212
rect 28320 -11268 28335 -11212
rect 28248 -11278 28335 -11268
rect 33095 -11212 33179 -11203
rect 33095 -11268 33111 -11212
rect 33167 -11268 33179 -11212
rect 33095 -11279 33179 -11268
rect 3665 -12107 3777 -12095
rect 3665 -12183 3688 -12107
rect 3758 -12183 3777 -12107
rect 3665 -12198 3777 -12183
rect 8523 -12114 8641 -12093
rect 8523 -12174 8559 -12114
rect 8617 -12174 8641 -12114
rect 8523 -12204 8641 -12174
rect 13474 -12116 13574 -12096
rect 13474 -12173 13504 -12116
rect 13564 -12173 13574 -12116
rect 13474 -12192 13574 -12173
rect 18221 -12118 18325 -12094
rect 18221 -12177 18249 -12118
rect 18313 -12177 18325 -12118
rect 18221 -12198 18325 -12177
rect 23150 -12113 23268 -12095
rect 23150 -12176 23190 -12113
rect 23255 -12176 23268 -12113
rect 23150 -12194 23268 -12176
rect 27977 -12117 28074 -12100
rect 27977 -12175 27998 -12117
rect 28058 -12175 28074 -12117
rect 27977 -12195 28074 -12175
rect 32865 -12116 32956 -12100
rect 32865 -12173 32888 -12116
rect 32944 -12173 32956 -12116
rect 32865 -12190 32956 -12173
rect 37731 -12114 37811 -12103
rect 37731 -12170 37744 -12114
rect 37800 -12170 37811 -12114
rect 37731 -12182 37811 -12170
rect 8391 -12589 8401 -12533
rect 8457 -12589 8467 -12533
rect 3453 -12880 3563 -12879
rect 8391 -12880 8467 -12589
rect 13240 -12585 13250 -12529
rect 13306 -12585 13316 -12529
rect 13240 -12880 13316 -12585
rect 18082 -12589 18092 -12533
rect 18148 -12589 18158 -12533
rect 18082 -12880 18158 -12589
rect 22922 -12593 22932 -12537
rect 22988 -12593 22998 -12537
rect 22922 -12880 22998 -12593
rect 27766 -12589 27776 -12533
rect 27832 -12589 27842 -12533
rect 27766 -12880 27842 -12589
rect 32638 -12592 32648 -12536
rect 32704 -12592 32714 -12536
rect 32638 -12880 32714 -12592
rect 37456 -12590 37466 -12534
rect 37522 -12590 37532 -12534
rect 37456 -12880 37532 -12590
rect 42662 -12712 42738 -12702
rect 42662 -12768 42672 -12712
rect 42728 -12768 42738 -12712
rect 42662 -12778 42738 -12768
rect 3136 -12940 39032 -12880
rect 3136 -12945 3469 -12940
rect 3136 -13001 3205 -12945
rect 3261 -12996 3469 -12945
rect 3525 -12996 4895 -12940
rect 4951 -12996 39032 -12940
rect 3261 -13001 39032 -12996
rect 3136 -13048 39032 -13001
rect 9762 -13340 9844 -13048
rect 9762 -13396 9774 -13340
rect 9830 -13396 9844 -13340
rect 14570 -13335 14655 -13048
rect 14570 -13391 14583 -13335
rect 14639 -13391 14655 -13335
rect 19448 -13333 19531 -13048
rect 19448 -13389 19461 -13333
rect 19517 -13389 19531 -13333
rect 24259 -13334 24344 -13048
rect 24259 -13390 24275 -13334
rect 24331 -13390 24344 -13334
rect 29135 -13332 29216 -13048
rect 29135 -13388 29148 -13332
rect 29204 -13388 29216 -13332
rect 33979 -13335 34061 -13048
rect 33979 -13391 33993 -13335
rect 34049 -13391 34061 -13335
rect 38823 -13335 38903 -13048
rect 38823 -13391 38837 -13335
rect 38893 -13391 38903 -13335
rect 4015 -14013 4108 -14001
rect 4015 -14070 4035 -14013
rect 4092 -14070 4108 -14013
rect 4015 -14078 4108 -14070
rect 8850 -14011 8968 -13998
rect 8850 -14069 8879 -14011
rect 8939 -14069 8968 -14011
rect 8850 -14080 8968 -14069
rect 13707 -14012 13799 -14005
rect 13707 -14069 13725 -14012
rect 13784 -14069 13799 -14012
rect 13707 -14079 13799 -14069
rect 18551 -14011 18649 -13996
rect 18551 -14068 18572 -14011
rect 18630 -14068 18649 -14011
rect 18551 -14088 18649 -14068
rect 23405 -14013 23488 -14001
rect 23405 -14070 23417 -14013
rect 23477 -14070 23488 -14013
rect 23405 -14080 23488 -14070
rect 28250 -14012 28333 -14003
rect 28250 -14068 28263 -14012
rect 28321 -14068 28333 -14012
rect 28250 -14076 28333 -14068
rect 33095 -14012 33178 -14005
rect 33095 -14069 33110 -14012
rect 33166 -14069 33178 -14012
rect 33095 -14078 33178 -14069
rect 3656 -14907 3771 -14898
rect 3656 -14983 3681 -14907
rect 3746 -14983 3771 -14907
rect 3656 -14995 3771 -14983
rect 8539 -14917 8649 -14896
rect 8539 -14973 8578 -14917
rect 8636 -14973 8649 -14917
rect 8539 -14997 8649 -14973
rect 13474 -14916 13578 -14897
rect 13474 -14973 13509 -14916
rect 13568 -14973 13578 -14916
rect 13474 -14991 13578 -14973
rect 18227 -14917 18340 -14891
rect 18227 -14979 18252 -14917
rect 18316 -14979 18340 -14917
rect 18227 -15005 18340 -14979
rect 23147 -14909 23265 -14892
rect 23147 -14974 23191 -14909
rect 23254 -14974 23265 -14909
rect 23147 -14996 23265 -14974
rect 27979 -14916 28076 -14899
rect 27979 -14972 27997 -14916
rect 28062 -14972 28076 -14916
rect 27979 -14989 28076 -14972
rect 32845 -14916 32949 -14904
rect 32845 -14974 32866 -14916
rect 32938 -14974 32949 -14916
rect 32845 -14989 32949 -14974
rect 37733 -14914 37812 -14903
rect 37733 -14970 37744 -14914
rect 37800 -14970 37812 -14914
rect 37733 -14981 37812 -14970
rect 27767 -15335 27843 -15334
rect 8392 -15393 8402 -15337
rect 8458 -15393 8468 -15337
rect 8392 -15680 8468 -15393
rect 13238 -15395 13248 -15339
rect 13304 -15395 13314 -15339
rect 13238 -15680 13314 -15395
rect 18081 -15391 18091 -15335
rect 18147 -15391 18157 -15335
rect 18081 -15680 18157 -15391
rect 22950 -15391 22960 -15335
rect 23016 -15391 23026 -15335
rect 22950 -15680 23026 -15391
rect 27767 -15391 27777 -15335
rect 27833 -15391 27843 -15335
rect 27767 -15680 27843 -15391
rect 32638 -15388 32648 -15332
rect 32704 -15388 32714 -15332
rect 32638 -15680 32714 -15388
rect 37454 -15387 37464 -15331
rect 37520 -15387 37530 -15331
rect 37454 -15680 37530 -15387
rect 42662 -15512 42738 -15502
rect 42662 -15568 42672 -15512
rect 42728 -15568 42738 -15512
rect 42662 -15578 42738 -15568
rect 3080 -15738 39032 -15680
rect 3080 -15794 3191 -15738
rect 3247 -15740 39032 -15738
rect 3247 -15746 4898 -15740
rect 3247 -15794 3471 -15746
rect 3080 -15802 3471 -15794
rect 3527 -15796 4898 -15746
rect 4954 -15796 39032 -15740
rect 3527 -15802 39032 -15796
rect 3080 -15848 39032 -15802
rect 9762 -16140 9844 -15848
rect 13238 -15849 13314 -15848
rect 9762 -16196 9774 -16140
rect 9830 -16196 9844 -16140
rect 14570 -16137 14655 -15848
rect 14570 -16193 14584 -16137
rect 14640 -16193 14655 -16137
rect 19448 -16135 19531 -15848
rect 19448 -16191 19463 -16135
rect 19519 -16191 19531 -16135
rect 24259 -16142 24344 -15848
rect 24259 -16198 24273 -16142
rect 24329 -16198 24344 -16142
rect 29135 -16134 29216 -15848
rect 29135 -16190 29148 -16134
rect 29204 -16190 29216 -16134
rect 33979 -16134 34061 -15848
rect 33979 -16190 33993 -16134
rect 34049 -16190 34061 -16134
rect 38823 -16135 38903 -15848
rect 38823 -16191 38835 -16135
rect 38891 -16191 38903 -16135
rect 4018 -16812 4107 -16806
rect 4018 -16868 4034 -16812
rect 4090 -16868 4107 -16812
rect 4018 -16876 4107 -16868
rect 8857 -16812 8959 -16805
rect 8857 -16870 8879 -16812
rect 8938 -16870 8959 -16812
rect 8857 -16879 8959 -16870
rect 13710 -16812 13795 -16806
rect 13710 -16869 13726 -16812
rect 13785 -16869 13795 -16812
rect 13710 -16881 13795 -16869
rect 18558 -16810 18643 -16799
rect 18558 -16869 18572 -16810
rect 18630 -16869 18643 -16810
rect 18558 -16884 18643 -16869
rect 23406 -16811 23491 -16801
rect 23406 -16870 23415 -16811
rect 23478 -16870 23491 -16811
rect 23406 -16880 23491 -16870
rect 28249 -16811 28334 -16804
rect 28249 -16867 28265 -16811
rect 28323 -16867 28334 -16811
rect 28249 -16875 28334 -16867
rect 33096 -16813 33184 -16801
rect 33096 -16870 33109 -16813
rect 33167 -16870 33184 -16813
rect 33096 -16878 33184 -16870
rect 3664 -17707 3776 -17696
rect 3664 -17783 3692 -17707
rect 3760 -17783 3776 -17707
rect 3664 -17796 3776 -17783
rect 8538 -17717 8646 -17693
rect 8538 -17775 8570 -17717
rect 8630 -17775 8646 -17717
rect 8538 -17798 8646 -17775
rect 13483 -17715 13572 -17699
rect 13483 -17771 13505 -17715
rect 13561 -17771 13572 -17715
rect 13483 -17793 13572 -17771
rect 18221 -17715 18335 -17695
rect 18221 -17776 18250 -17715
rect 18318 -17776 18335 -17715
rect 18221 -17796 18335 -17776
rect 23153 -17712 23267 -17694
rect 23153 -17778 23191 -17712
rect 23251 -17778 23267 -17712
rect 23153 -17798 23267 -17778
rect 27983 -17712 28077 -17698
rect 27983 -17769 27999 -17712
rect 28060 -17769 28077 -17712
rect 27983 -17787 28077 -17769
rect 32850 -17715 32945 -17702
rect 32850 -17775 32868 -17715
rect 32935 -17775 32945 -17715
rect 32850 -17791 32945 -17775
rect 37735 -17716 37813 -17703
rect 37735 -17772 37744 -17716
rect 37800 -17772 37813 -17716
rect 37735 -17783 37813 -17772
rect 8390 -18193 8400 -18137
rect 8456 -18193 8466 -18137
rect 8390 -18480 8466 -18193
rect 13252 -18196 13262 -18140
rect 13318 -18196 13328 -18140
rect 13252 -18480 13328 -18196
rect 18080 -18190 18090 -18134
rect 18146 -18190 18156 -18134
rect 18080 -18480 18156 -18190
rect 22946 -18190 22956 -18134
rect 23012 -18190 23022 -18134
rect 22946 -18480 23022 -18190
rect 27769 -18192 27779 -18136
rect 27835 -18192 27845 -18136
rect 27769 -18480 27845 -18192
rect 32636 -18194 32646 -18138
rect 32702 -18194 32712 -18138
rect 32636 -18480 32712 -18194
rect 37456 -18480 37532 -18197
rect 42662 -18312 42738 -18302
rect 42662 -18368 42672 -18312
rect 42728 -18368 42738 -18312
rect 42662 -18378 42738 -18368
rect 3416 -18513 39032 -18480
rect 3416 -18569 3471 -18513
rect 3527 -18569 39032 -18513
rect 3416 -18648 39032 -18569
rect 4883 -19499 4966 -18648
rect 4883 -19555 4893 -19499
rect 4956 -19555 4966 -19499
rect 4883 -19561 4966 -19555
rect 9762 -19498 9844 -18648
rect 9762 -19554 9772 -19498
rect 9834 -19554 9844 -19498
rect 9762 -19561 9844 -19554
rect 14570 -19501 14655 -18648
rect 14570 -19557 14580 -19501
rect 14645 -19557 14655 -19501
rect 14570 -19561 14655 -19557
rect 19448 -19502 19531 -18648
rect 19448 -19558 19458 -19502
rect 19521 -19558 19531 -19502
rect 19448 -19561 19531 -19558
rect 24259 -19499 24344 -18648
rect 24259 -19556 24269 -19499
rect 24334 -19556 24344 -19499
rect 24259 -19561 24344 -19556
rect 29135 -19502 29216 -18648
rect 29135 -19558 29145 -19502
rect 29206 -19558 29216 -19502
rect 33979 -19501 34061 -18648
rect 37456 -18649 37532 -18648
rect 38823 -18649 38903 -18648
rect 33979 -19557 33989 -19501
rect 34051 -19557 34061 -19501
rect 33979 -19561 34061 -19557
rect 4018 -19613 4107 -19608
rect 4018 -19669 4034 -19613
rect 4091 -19669 4107 -19613
rect 4018 -19678 4107 -19669
rect 8862 -19612 8956 -19603
rect 8862 -19668 8881 -19612
rect 8939 -19668 8956 -19612
rect 8862 -19678 8956 -19668
rect 13713 -19612 13794 -19602
rect 13713 -19668 13727 -19612
rect 13784 -19668 13794 -19612
rect 13713 -19676 13794 -19668
rect 18555 -19613 18649 -19595
rect 18555 -19669 18573 -19613
rect 18630 -19669 18649 -19613
rect 18555 -19683 18649 -19669
rect 23404 -19612 23485 -19605
rect 23404 -19669 23417 -19612
rect 23476 -19669 23485 -19612
rect 23404 -19679 23485 -19669
rect 28246 -19612 28338 -19599
rect 28246 -19669 28262 -19612
rect 28319 -19669 28338 -19612
rect 28246 -19681 28338 -19669
rect 33090 -19611 33189 -19600
rect 33090 -19670 33108 -19611
rect 33170 -19670 33189 -19611
rect 33090 -19685 33189 -19670
rect 3664 -20507 3772 -20496
rect 3664 -20583 3696 -20507
rect 3752 -20583 3772 -20507
rect 3664 -20596 3772 -20583
rect 8532 -20514 8651 -20494
rect 8532 -20573 8563 -20514
rect 8625 -20573 8651 -20514
rect 8532 -20601 8651 -20573
rect 13484 -20515 13581 -20501
rect 13484 -20571 13513 -20515
rect 13571 -20571 13581 -20515
rect 13484 -20589 13581 -20571
rect 18223 -20518 18334 -20497
rect 18223 -20580 18251 -20518
rect 18315 -20580 18334 -20518
rect 18223 -20598 18334 -20580
rect 23162 -20514 23270 -20496
rect 23162 -20577 23193 -20514
rect 23253 -20577 23270 -20514
rect 23162 -20597 23270 -20577
rect 27983 -20517 28072 -20496
rect 27983 -20574 27998 -20517
rect 28059 -20574 28072 -20517
rect 27983 -20587 28072 -20574
rect 32859 -20517 32943 -20503
rect 32859 -20574 32869 -20517
rect 32932 -20574 32943 -20517
rect 32859 -20586 32943 -20574
rect 42662 -21112 42738 -21102
rect 42662 -21168 42672 -21112
rect 42728 -21168 42738 -21112
rect 42662 -21178 42738 -21168
<< via3 >>
rect 3696 2436 3752 2492
rect 8568 2436 8624 2492
rect 13496 2438 13552 2494
rect 18256 2435 18312 2491
rect 23184 2436 23240 2492
rect 28000 2441 28056 2497
rect 32872 2408 32928 2464
rect 37744 2408 37800 2464
rect 13716 1203 13780 1278
rect 18562 1185 18631 1257
rect 23403 1223 23468 1301
rect 28271 1218 28344 1291
rect 33095 1202 33156 1262
rect 8856 813 8928 876
rect 4029 480 4093 537
rect 4033 -69 4092 -13
rect 8880 -68 8938 -12
rect 13725 -69 13784 -13
rect 18570 -70 18632 -12
rect 23418 -69 23476 -12
rect 28262 -69 28325 -13
rect 33109 -70 33168 -13
rect 3696 -983 3774 -907
rect 8574 -983 8632 -907
rect 13505 -974 13567 -916
rect 18256 -972 18315 -915
rect 23194 -971 23260 -913
rect 27999 -975 28058 -915
rect 32869 -972 32932 -915
rect 37744 -971 37800 -915
rect 42672 -1568 42728 -1512
rect 4035 -2868 4092 -2812
rect 8879 -2870 8938 -2812
rect 13725 -2869 13784 -2812
rect 18570 -2870 18629 -2812
rect 23416 -2870 23475 -2813
rect 28265 -2868 28322 -2810
rect 33110 -2869 33166 -2813
rect 3687 -3783 3755 -3707
rect 8568 -3783 8628 -3707
rect 13507 -3774 13570 -3714
rect 18259 -3777 18323 -3716
rect 23194 -3774 23253 -3718
rect 27990 -3772 28052 -3714
rect 32869 -3774 32932 -3714
rect 37744 -3770 37800 -3714
rect 42672 -4368 42728 -4312
rect 4035 -5668 4091 -5612
rect 8878 -5670 8937 -5613
rect 13725 -5669 13783 -5613
rect 18569 -5671 18634 -5607
rect 23416 -5671 23478 -5610
rect 28264 -5668 28323 -5611
rect 33109 -5669 33169 -5611
rect 3691 -6583 3750 -6507
rect 8565 -6583 8624 -6507
rect 13506 -6573 13569 -6513
rect 18253 -6577 18318 -6517
rect 23194 -6572 23252 -6516
rect 27985 -6576 28045 -6515
rect 32870 -6573 32933 -6517
rect 37744 -6570 37800 -6514
rect 42671 -7168 42728 -7112
rect 4034 -8469 4091 -8413
rect 8878 -8471 8942 -8411
rect 13726 -8469 13782 -8413
rect 18571 -8470 18629 -8412
rect 23416 -8471 23479 -8406
rect 28262 -8469 28323 -8411
rect 33107 -8471 33166 -8413
rect 3696 -9373 3752 -9317
rect 8566 -9383 8627 -9307
rect 13505 -9373 13570 -9314
rect 18252 -9376 18318 -9317
rect 23194 -9373 23252 -9314
rect 27993 -9375 28053 -9317
rect 32867 -9374 32933 -9316
rect 37744 -9371 37800 -9315
rect 42672 -9968 42728 -9912
rect 4035 -11268 4091 -11212
rect 8874 -11272 8938 -11212
rect 13726 -11269 13782 -11212
rect 18571 -11270 18630 -11210
rect 23417 -11270 23480 -11210
rect 28264 -11268 28320 -11212
rect 33111 -11268 33167 -11212
rect 3688 -12183 3758 -12107
rect 8559 -12174 8617 -12114
rect 13504 -12173 13564 -12116
rect 18249 -12177 18313 -12118
rect 23190 -12176 23255 -12113
rect 27998 -12175 28058 -12117
rect 32888 -12173 32944 -12116
rect 37744 -12170 37800 -12114
rect 42672 -12768 42728 -12712
rect 4035 -14070 4092 -14013
rect 8879 -14069 8939 -14011
rect 13725 -14069 13784 -14012
rect 18572 -14068 18630 -14011
rect 23417 -14070 23477 -14013
rect 28263 -14068 28321 -14012
rect 33110 -14069 33166 -14012
rect 3681 -14983 3746 -14907
rect 8578 -14973 8636 -14917
rect 13509 -14973 13568 -14916
rect 18252 -14979 18316 -14917
rect 23191 -14974 23254 -14909
rect 27997 -14972 28062 -14916
rect 32866 -14974 32938 -14916
rect 37744 -14970 37800 -14914
rect 42672 -15568 42728 -15512
rect 4034 -16868 4090 -16812
rect 8879 -16870 8938 -16812
rect 13726 -16869 13785 -16812
rect 18572 -16869 18630 -16810
rect 23415 -16870 23478 -16811
rect 28265 -16867 28323 -16811
rect 33109 -16870 33167 -16813
rect 3692 -17783 3760 -17707
rect 8570 -17775 8630 -17717
rect 13505 -17771 13561 -17715
rect 18250 -17776 18318 -17715
rect 23191 -17778 23251 -17712
rect 27999 -17769 28060 -17712
rect 32868 -17775 32935 -17715
rect 37744 -17772 37800 -17716
rect 42672 -18368 42728 -18312
rect 4034 -19669 4091 -19613
rect 8881 -19668 8939 -19612
rect 13727 -19668 13784 -19612
rect 18573 -19669 18630 -19613
rect 23417 -19669 23476 -19612
rect 28262 -19669 28319 -19612
rect 33108 -19670 33170 -19611
rect 3696 -20583 3752 -20507
rect 8563 -20573 8625 -20514
rect 13513 -20571 13571 -20515
rect 18251 -20580 18315 -20518
rect 23193 -20577 23253 -20514
rect 27998 -20574 28059 -20517
rect 32869 -20574 32932 -20517
rect 42672 -21168 42728 -21112
<< metal4 >>
rect 3640 2492 3808 2632
rect 3640 2436 3696 2492
rect 3752 2436 3808 2492
rect 3640 -907 3808 2436
rect 8512 2492 8680 2632
rect 8512 2436 8568 2492
rect 8624 2436 8680 2492
rect 3640 -983 3696 -907
rect 3774 -983 3808 -907
rect 3640 -3707 3808 -983
rect 3640 -3783 3687 -3707
rect 3755 -3783 3808 -3707
rect 3640 -6507 3808 -3783
rect 3640 -6583 3691 -6507
rect 3750 -6583 3808 -6507
rect 3640 -9317 3808 -6583
rect 3640 -9373 3696 -9317
rect 3752 -9373 3808 -9317
rect 3640 -12107 3808 -9373
rect 3640 -12183 3688 -12107
rect 3758 -12183 3808 -12107
rect 3640 -14907 3808 -12183
rect 3640 -14983 3681 -14907
rect 3746 -14983 3808 -14907
rect 3640 -17707 3808 -14983
rect 3640 -17783 3692 -17707
rect 3760 -17783 3808 -17707
rect 3640 -20507 3808 -17783
rect 3640 -20583 3696 -20507
rect 3752 -20583 3808 -20507
rect 3640 -21224 3808 -20583
rect 3976 537 4144 560
rect 3976 480 4029 537
rect 4093 480 4144 537
rect 3976 -13 4144 480
rect 3976 -69 4033 -13
rect 4092 -69 4144 -13
rect 3976 -2812 4144 -69
rect 3976 -2868 4035 -2812
rect 4092 -2868 4144 -2812
rect 3976 -5612 4144 -2868
rect 3976 -5668 4035 -5612
rect 4091 -5668 4144 -5612
rect 3976 -8413 4144 -5668
rect 3976 -8469 4034 -8413
rect 4091 -8469 4144 -8413
rect 3976 -11212 4144 -8469
rect 3976 -11268 4035 -11212
rect 4091 -11268 4144 -11212
rect 3976 -14013 4144 -11268
rect 3976 -14070 4035 -14013
rect 4092 -14070 4144 -14013
rect 3976 -16812 4144 -14070
rect 3976 -16868 4034 -16812
rect 4090 -16868 4144 -16812
rect 3976 -19613 4144 -16868
rect 3976 -19669 4034 -19613
rect 4091 -19669 4144 -19613
rect 3976 -21224 4144 -19669
rect 8512 -907 8680 2436
rect 13440 2494 13608 2632
rect 13440 2438 13496 2494
rect 13552 2438 13608 2494
rect 8512 -983 8574 -907
rect 8632 -983 8680 -907
rect 8512 -3707 8680 -983
rect 8512 -3783 8568 -3707
rect 8628 -3783 8680 -3707
rect 8512 -6507 8680 -3783
rect 8512 -6583 8565 -6507
rect 8624 -6583 8680 -6507
rect 8512 -9307 8680 -6583
rect 8512 -9383 8566 -9307
rect 8627 -9383 8680 -9307
rect 8512 -12114 8680 -9383
rect 8512 -12174 8559 -12114
rect 8617 -12174 8680 -12114
rect 8512 -14917 8680 -12174
rect 8512 -14973 8578 -14917
rect 8636 -14973 8680 -14917
rect 8512 -17717 8680 -14973
rect 8512 -17775 8570 -17717
rect 8630 -17775 8680 -17717
rect 8512 -20514 8680 -17775
rect 8512 -20573 8563 -20514
rect 8625 -20573 8680 -20514
rect 8512 -21392 8680 -20573
rect 8818 876 8996 1039
rect 8818 813 8856 876
rect 8928 813 8996 876
rect 8818 -12 8996 813
rect 8818 -68 8880 -12
rect 8938 -68 8996 -12
rect 8818 -2812 8996 -68
rect 8818 -2870 8879 -2812
rect 8938 -2870 8996 -2812
rect 8818 -5613 8996 -2870
rect 8818 -5670 8878 -5613
rect 8937 -5670 8996 -5613
rect 8818 -8411 8996 -5670
rect 8818 -8471 8878 -8411
rect 8942 -8471 8996 -8411
rect 8818 -11212 8996 -8471
rect 8818 -11272 8874 -11212
rect 8938 -11272 8996 -11212
rect 8818 -14011 8996 -11272
rect 8818 -14069 8879 -14011
rect 8939 -14069 8996 -14011
rect 8818 -16812 8996 -14069
rect 8818 -16870 8879 -16812
rect 8938 -16870 8996 -16812
rect 8818 -19612 8996 -16870
rect 8818 -19668 8881 -19612
rect 8939 -19668 8996 -19612
rect 8818 -21392 8996 -19668
rect 13440 -916 13608 2438
rect 18200 2491 18368 2632
rect 18200 2435 18256 2491
rect 18312 2435 18368 2491
rect 13440 -974 13505 -916
rect 13567 -974 13608 -916
rect 13440 -3714 13608 -974
rect 13440 -3774 13507 -3714
rect 13570 -3774 13608 -3714
rect 13440 -6513 13608 -3774
rect 13440 -6573 13506 -6513
rect 13569 -6573 13608 -6513
rect 13440 -9314 13608 -6573
rect 13440 -9373 13505 -9314
rect 13570 -9373 13608 -9314
rect 13440 -12116 13608 -9373
rect 13440 -12173 13504 -12116
rect 13564 -12173 13608 -12116
rect 13440 -14916 13608 -12173
rect 13440 -14973 13509 -14916
rect 13568 -14973 13608 -14916
rect 13440 -17715 13608 -14973
rect 13440 -17771 13505 -17715
rect 13561 -17771 13608 -17715
rect 13440 -20515 13608 -17771
rect 13440 -20571 13513 -20515
rect 13571 -20571 13608 -20515
rect 13440 -21336 13608 -20571
rect 13664 1278 13832 1344
rect 13664 1203 13716 1278
rect 13780 1203 13832 1278
rect 13664 952 13832 1203
rect 13664 -13 13833 952
rect 13664 -69 13725 -13
rect 13784 -69 13833 -13
rect 13664 -2812 13833 -69
rect 13664 -2869 13725 -2812
rect 13784 -2869 13833 -2812
rect 13664 -5613 13833 -2869
rect 13664 -5669 13725 -5613
rect 13783 -5669 13833 -5613
rect 13664 -8413 13833 -5669
rect 13664 -8469 13726 -8413
rect 13782 -8469 13833 -8413
rect 13664 -11212 13833 -8469
rect 13664 -11269 13726 -11212
rect 13782 -11269 13833 -11212
rect 13664 -14012 13833 -11269
rect 13664 -14069 13725 -14012
rect 13784 -14069 13833 -14012
rect 13664 -16812 13833 -14069
rect 13664 -16869 13726 -16812
rect 13785 -16869 13833 -16812
rect 13664 -19612 13833 -16869
rect 13664 -19668 13727 -19612
rect 13784 -19668 13833 -19612
rect 13664 -21336 13833 -19668
rect 18200 -915 18368 2435
rect 23128 2492 23296 2632
rect 23128 2436 23184 2492
rect 23240 2436 23296 2492
rect 18200 -972 18256 -915
rect 18315 -972 18368 -915
rect 18200 -3716 18368 -972
rect 18200 -3777 18259 -3716
rect 18323 -3777 18368 -3716
rect 18200 -6517 18368 -3777
rect 18200 -6577 18253 -6517
rect 18318 -6577 18368 -6517
rect 18200 -9317 18368 -6577
rect 18200 -9376 18252 -9317
rect 18318 -9376 18368 -9317
rect 18200 -12118 18368 -9376
rect 18200 -12177 18249 -12118
rect 18313 -12177 18368 -12118
rect 18200 -14917 18368 -12177
rect 18200 -14979 18252 -14917
rect 18316 -14979 18368 -14917
rect 18200 -17715 18368 -14979
rect 18200 -17776 18250 -17715
rect 18318 -17776 18368 -17715
rect 18200 -20518 18368 -17776
rect 18200 -20580 18251 -20518
rect 18315 -20580 18368 -20518
rect 18200 -21336 18368 -20580
rect 18505 1257 18674 1278
rect 18505 1185 18562 1257
rect 18631 1185 18674 1257
rect 18505 -12 18674 1185
rect 18505 -70 18570 -12
rect 18632 -70 18674 -12
rect 18505 -2812 18674 -70
rect 18505 -2870 18570 -2812
rect 18629 -2870 18674 -2812
rect 18505 -5607 18674 -2870
rect 18505 -5671 18569 -5607
rect 18634 -5671 18674 -5607
rect 18505 -8412 18674 -5671
rect 18505 -8470 18571 -8412
rect 18629 -8470 18674 -8412
rect 18505 -11210 18674 -8470
rect 18505 -11270 18571 -11210
rect 18630 -11270 18674 -11210
rect 18505 -14011 18674 -11270
rect 18505 -14068 18572 -14011
rect 18630 -14068 18674 -14011
rect 18505 -16810 18674 -14068
rect 18505 -16869 18572 -16810
rect 18630 -16869 18674 -16810
rect 18505 -19613 18674 -16869
rect 18505 -19669 18573 -19613
rect 18630 -19669 18674 -19613
rect 18505 -21336 18674 -19669
rect 23128 -913 23296 2436
rect 27944 2497 28112 2632
rect 27944 2441 28000 2497
rect 28056 2441 28112 2497
rect 23128 -971 23194 -913
rect 23260 -971 23296 -913
rect 23128 -3718 23296 -971
rect 23128 -3774 23194 -3718
rect 23253 -3774 23296 -3718
rect 23128 -6516 23296 -3774
rect 23128 -6572 23194 -6516
rect 23252 -6572 23296 -6516
rect 23128 -9314 23296 -6572
rect 23128 -9373 23194 -9314
rect 23252 -9373 23296 -9314
rect 23128 -12113 23296 -9373
rect 23128 -12176 23190 -12113
rect 23255 -12176 23296 -12113
rect 23128 -14909 23296 -12176
rect 23128 -14974 23191 -14909
rect 23254 -14974 23296 -14909
rect 23128 -17712 23296 -14974
rect 23128 -17778 23191 -17712
rect 23251 -17778 23296 -17712
rect 23128 -20514 23296 -17778
rect 23128 -20577 23193 -20514
rect 23253 -20577 23296 -20514
rect 23128 -21336 23296 -20577
rect 23352 1301 23520 1344
rect 23352 1223 23403 1301
rect 23468 1223 23520 1301
rect 23352 -12 23520 1223
rect 23352 -69 23418 -12
rect 23476 -69 23520 -12
rect 23352 -2813 23520 -69
rect 23352 -2870 23416 -2813
rect 23475 -2870 23520 -2813
rect 23352 -5610 23520 -2870
rect 23352 -5671 23416 -5610
rect 23478 -5671 23520 -5610
rect 23352 -8406 23520 -5671
rect 23352 -8471 23416 -8406
rect 23479 -8471 23520 -8406
rect 23352 -11210 23520 -8471
rect 23352 -11270 23417 -11210
rect 23480 -11270 23520 -11210
rect 23352 -14013 23520 -11270
rect 23352 -14070 23417 -14013
rect 23477 -14070 23520 -14013
rect 23352 -16811 23520 -14070
rect 23352 -16870 23415 -16811
rect 23478 -16870 23520 -16811
rect 23352 -19612 23520 -16870
rect 23352 -19669 23417 -19612
rect 23476 -19669 23520 -19612
rect 23352 -21336 23520 -19669
rect 27944 -915 28112 2441
rect 32816 2464 32984 2632
rect 32816 2408 32872 2464
rect 32928 2408 32984 2464
rect 27944 -975 27999 -915
rect 28058 -975 28112 -915
rect 27944 -3714 28112 -975
rect 27944 -3772 27990 -3714
rect 28052 -3772 28112 -3714
rect 27944 -6515 28112 -3772
rect 27944 -6576 27985 -6515
rect 28045 -6576 28112 -6515
rect 27944 -9317 28112 -6576
rect 27944 -9375 27993 -9317
rect 28053 -9375 28112 -9317
rect 27944 -12117 28112 -9375
rect 27944 -12175 27998 -12117
rect 28058 -12175 28112 -12117
rect 27944 -14916 28112 -12175
rect 27944 -14972 27997 -14916
rect 28062 -14972 28112 -14916
rect 27944 -17712 28112 -14972
rect 27944 -17769 27999 -17712
rect 28060 -17769 28112 -17712
rect 27944 -20517 28112 -17769
rect 27944 -20574 27998 -20517
rect 28059 -20574 28112 -20517
rect 27944 -21336 28112 -20574
rect 28224 1291 28392 1336
rect 28224 1218 28271 1291
rect 28344 1218 28392 1291
rect 28224 -13 28392 1218
rect 28224 -69 28262 -13
rect 28325 -69 28392 -13
rect 28224 -2810 28392 -69
rect 28224 -2868 28265 -2810
rect 28322 -2868 28392 -2810
rect 28224 -5611 28392 -2868
rect 28224 -5668 28264 -5611
rect 28323 -5668 28392 -5611
rect 28224 -8411 28392 -5668
rect 28224 -8469 28262 -8411
rect 28323 -8469 28392 -8411
rect 28224 -11212 28392 -8469
rect 28224 -11268 28264 -11212
rect 28320 -11268 28392 -11212
rect 28224 -14012 28392 -11268
rect 28224 -14068 28263 -14012
rect 28321 -14068 28392 -14012
rect 28224 -16811 28392 -14068
rect 28224 -16867 28265 -16811
rect 28323 -16867 28392 -16811
rect 28224 -19612 28392 -16867
rect 28224 -19669 28262 -19612
rect 28319 -19669 28392 -19612
rect 28224 -21336 28392 -19669
rect 32816 -915 32984 2408
rect 37688 2464 37856 2576
rect 37688 2408 37744 2464
rect 37800 2408 37856 2464
rect 32816 -972 32869 -915
rect 32932 -972 32984 -915
rect 32816 -3714 32984 -972
rect 32816 -3774 32869 -3714
rect 32932 -3774 32984 -3714
rect 32816 -6517 32984 -3774
rect 32816 -6573 32870 -6517
rect 32933 -6573 32984 -6517
rect 32816 -9316 32984 -6573
rect 32816 -9374 32867 -9316
rect 32933 -9374 32984 -9316
rect 32816 -12116 32984 -9374
rect 32816 -12173 32888 -12116
rect 32944 -12173 32984 -12116
rect 32816 -14916 32984 -12173
rect 32816 -14974 32866 -14916
rect 32938 -14974 32984 -14916
rect 32816 -17715 32984 -14974
rect 32816 -17775 32868 -17715
rect 32935 -17775 32984 -17715
rect 32816 -20517 32984 -17775
rect 32816 -20574 32869 -20517
rect 32932 -20574 32984 -20517
rect 32816 -21392 32984 -20574
rect 33040 1262 33208 1288
rect 33040 1202 33095 1262
rect 33156 1202 33208 1262
rect 33040 -13 33208 1202
rect 33040 -70 33109 -13
rect 33168 -70 33208 -13
rect 33040 -2813 33208 -70
rect 33040 -2869 33110 -2813
rect 33166 -2869 33208 -2813
rect 33040 -5611 33208 -2869
rect 33040 -5669 33109 -5611
rect 33169 -5669 33208 -5611
rect 33040 -8413 33208 -5669
rect 33040 -8471 33107 -8413
rect 33166 -8471 33208 -8413
rect 33040 -11212 33208 -8471
rect 33040 -11268 33111 -11212
rect 33167 -11268 33208 -11212
rect 33040 -14012 33208 -11268
rect 33040 -14069 33110 -14012
rect 33166 -14069 33208 -14012
rect 33040 -16813 33208 -14069
rect 33040 -16870 33109 -16813
rect 33167 -16870 33208 -16813
rect 33040 -19611 33208 -16870
rect 37688 -915 37856 2408
rect 37688 -971 37744 -915
rect 37800 -971 37856 -915
rect 37688 -3714 37856 -971
rect 37688 -3770 37744 -3714
rect 37800 -3770 37856 -3714
rect 37688 -6514 37856 -3770
rect 37688 -6570 37744 -6514
rect 37800 -6570 37856 -6514
rect 37688 -9315 37856 -6570
rect 37688 -9371 37744 -9315
rect 37800 -9371 37856 -9315
rect 37688 -12114 37856 -9371
rect 37688 -12170 37744 -12114
rect 37800 -12170 37856 -12114
rect 37688 -14914 37856 -12170
rect 37688 -14970 37744 -14914
rect 37800 -14970 37856 -14914
rect 37688 -17716 37856 -14970
rect 37688 -17772 37744 -17716
rect 37800 -17772 37856 -17716
rect 37688 -18032 37856 -17772
rect 42560 -1512 42896 1400
rect 42560 -1568 42672 -1512
rect 42728 -1568 42896 -1512
rect 42560 -4312 42896 -1568
rect 42560 -4368 42672 -4312
rect 42728 -4368 42896 -4312
rect 42560 -7112 42896 -4368
rect 42560 -7168 42671 -7112
rect 42728 -7168 42896 -7112
rect 42560 -9912 42896 -7168
rect 42560 -9968 42672 -9912
rect 42728 -9968 42896 -9912
rect 42560 -12712 42896 -9968
rect 42560 -12768 42672 -12712
rect 42728 -12768 42896 -12712
rect 42560 -15512 42896 -12768
rect 42560 -15568 42672 -15512
rect 42728 -15568 42896 -15512
rect 33040 -19670 33108 -19611
rect 33170 -19670 33208 -19611
rect 33040 -21392 33208 -19670
rect 42560 -18312 42896 -15568
rect 42560 -18368 42672 -18312
rect 42728 -18368 42896 -18312
rect 42560 -21112 42896 -18368
rect 42560 -21168 42672 -21112
rect 42728 -21168 42896 -21112
rect 42560 -21392 42896 -21168
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2506 0 1 -12537
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_1
timestamp 1753044640
transform 1 0 2384 0 -1 -5249
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_2
timestamp 1753044640
transform 1 0 2490 0 1 -18137
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_3
timestamp 1753044640
transform 1 0 2493 0 1 -15337
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_4
timestamp 1753044640
transform 1 0 2490 0 -1 -16449
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_5
timestamp 1753044640
transform 1 0 22038 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_6
timestamp 1753044640
transform 1 0 11286 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_7
timestamp 1753044640
transform 1 0 27078 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_8
timestamp 1753044640
transform 1 0 31726 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  gf180mcu_fd_sc_mcu7t5v0__and2_2_9
timestamp 1753044640
transform 1 0 30606 0 1 1038
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2602 0 1 -9737
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  gf180mcu_fd_sc_mcu7t5v0__buf_2_1
timestamp 1753044640
transform 1 0 17278 0 1 1038
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_0 ~/eda/unic-cass/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2403 0 -1 351
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_1
timestamp 1753044640
transform 1 0 2388 0 1 -4137
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_2
timestamp 1753044640
transform 1 0 2403 0 1 -1337
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_3
timestamp 1753044640
transform 1 0 2394 0 -1 -10849
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_4
timestamp 1753044640
transform 1 0 2384 0 1 -6937
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_5
timestamp 1753044640
transform 1 0 2403 0 1 471
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_6
timestamp 1753044640
transform 1 0 2403 0 -1 2159
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_7
timestamp 1753044640
transform 1 0 6022 0 1 471
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_8
timestamp 1753044640
transform 1 0 20918 0 1 1038
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  gf180mcu_fd_sc_mcu7t5v0__or2_2_9
timestamp 1753044640
transform 1 0 12294 0 1 1038
box -86 -86 1206 870
use unit_cell_array  unit_cell_array_0
timestamp 1755843645
transform 1 0 13288 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_1
timestamp 1755843645
transform 1 0 3596 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_2
timestamp 1755843645
transform 1 0 8442 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_3
timestamp 1755843645
transform 1 0 37518 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_4
timestamp 1755843645
transform 1 0 18134 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_5
timestamp 1755843645
transform 1 0 22980 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_6
timestamp 1755843645
transform 1 0 27826 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_7
timestamp 1755843645
transform 1 0 32672 0 1 -254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_8
timestamp 1755843645
transform 1 0 8442 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_9
timestamp 1755843645
transform 1 0 3596 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_10
timestamp 1755843645
transform 1 0 13288 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_11
timestamp 1755843645
transform 1 0 22980 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_12
timestamp 1755843645
transform 1 0 18134 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_13
timestamp 1755843645
transform 1 0 27826 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_14
timestamp 1755843645
transform 1 0 37518 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_15
timestamp 1755843645
transform 1 0 32672 0 1 -3054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_17
timestamp 1755843645
transform 1 0 32672 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_18
timestamp 1755843645
transform 1 0 27826 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_19
timestamp 1755843645
transform 1 0 22980 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_20
timestamp 1755843645
transform 1 0 18134 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_21
timestamp 1755843645
transform 1 0 13288 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_22
timestamp 1755843645
transform 1 0 8442 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_23
timestamp 1755843645
transform 1 0 3596 0 1 -19854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_24
timestamp 1755843645
transform 1 0 8442 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_25
timestamp 1755843645
transform 1 0 3596 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_26
timestamp 1755843645
transform 1 0 13288 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_27
timestamp 1755843645
transform 1 0 22980 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_28
timestamp 1755843645
transform 1 0 18134 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_29
timestamp 1755843645
transform 1 0 27826 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_30
timestamp 1755843645
transform 1 0 37518 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_31
timestamp 1755843645
transform 1 0 32672 0 1 -5854
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_32
timestamp 1755843645
transform 1 0 8442 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_33
timestamp 1755843645
transform 1 0 3596 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_34
timestamp 1755843645
transform 1 0 13288 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_35
timestamp 1755843645
transform 1 0 22980 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_36
timestamp 1755843645
transform 1 0 18134 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_37
timestamp 1755843645
transform 1 0 27826 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_38
timestamp 1755843645
transform 1 0 37518 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_39
timestamp 1755843645
transform 1 0 32672 0 1 -8654
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_40
timestamp 1755843645
transform 1 0 8442 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_41
timestamp 1755843645
transform 1 0 3596 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_42
timestamp 1755843645
transform 1 0 13288 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_43
timestamp 1755843645
transform 1 0 22980 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_44
timestamp 1755843645
transform 1 0 18134 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_45
timestamp 1755843645
transform 1 0 27826 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_46
timestamp 1755843645
transform 1 0 37518 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_47
timestamp 1755843645
transform 1 0 32672 0 1 -11454
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_48
timestamp 1755843645
transform 1 0 8442 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_49
timestamp 1755843645
transform 1 0 3596 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_50
timestamp 1755843645
transform 1 0 13288 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_51
timestamp 1755843645
transform 1 0 22980 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_52
timestamp 1755843645
transform 1 0 18134 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_53
timestamp 1755843645
transform 1 0 27826 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_54
timestamp 1755843645
transform 1 0 37518 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_55
timestamp 1755843645
transform 1 0 32672 0 1 -14254
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_56
timestamp 1755843645
transform 1 0 8442 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_57
timestamp 1755843645
transform 1 0 3596 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_58
timestamp 1755843645
transform 1 0 13288 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_59
timestamp 1755843645
transform 1 0 22980 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_60
timestamp 1755843645
transform 1 0 18134 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_61
timestamp 1755843645
transform 1 0 27826 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_62
timestamp 1755843645
transform 1 0 37518 0 1 -17054
box -12 -1202 4834 691
use unit_cell_array  unit_cell_array_63
timestamp 1755843645
transform 1 0 32672 0 1 -17054
box -12 -1202 4834 691
<< end >>
