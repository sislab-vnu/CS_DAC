magic
tech gf180mcuD
magscale 1 10
timestamp 1754379792
<< pwell >>
rect -326 -1889 1387 -1024
<< nmos >>
rect -56 -1512 0 -1468
rect 172 -1511 228 -1467
rect 557 -1507 613 -1463
rect 705 -1507 1145 -1463
<< ndiff >>
rect -181 -1465 -101 -1448
rect -181 -1512 -164 -1465
rect -118 -1468 -101 -1465
rect 46 -1465 126 -1448
rect 46 -1468 63 -1465
rect -118 -1512 -56 -1468
rect 0 -1512 63 -1468
rect 109 -1467 126 -1465
rect 273 -1467 353 -1451
rect 109 -1511 172 -1467
rect 228 -1468 353 -1467
rect 228 -1511 290 -1468
rect 109 -1512 126 -1511
rect -181 -1529 -101 -1512
rect 46 -1529 126 -1512
rect 273 -1515 290 -1511
rect 336 -1515 353 -1468
rect 273 -1532 353 -1515
rect 432 -1462 512 -1445
rect 432 -1509 449 -1462
rect 495 -1463 512 -1462
rect 1191 -1462 1271 -1445
rect 1191 -1463 1208 -1462
rect 495 -1507 557 -1463
rect 613 -1507 705 -1463
rect 1145 -1507 1208 -1463
rect 495 -1509 512 -1507
rect 432 -1526 512 -1509
rect 1191 -1509 1208 -1507
rect 1254 -1509 1271 -1462
rect 1191 -1526 1271 -1509
<< ndiffc >>
rect -164 -1512 -118 -1465
rect 63 -1512 109 -1465
rect 290 -1515 336 -1468
rect 449 -1509 495 -1462
rect 1208 -1509 1254 -1462
<< polysilicon >>
rect -70 -1361 10 -1341
rect -70 -1408 -52 -1361
rect -6 -1408 10 -1361
rect -70 -1422 10 -1408
rect 160 -1361 240 -1341
rect 160 -1408 178 -1361
rect 224 -1408 240 -1361
rect 160 -1422 240 -1408
rect 557 -1384 1144 -1343
rect -56 -1468 0 -1422
rect 172 -1467 228 -1422
rect 557 -1424 865 -1384
rect -56 -1558 0 -1512
rect 172 -1557 228 -1511
rect 557 -1463 613 -1424
rect 705 -1430 865 -1424
rect 985 -1417 1144 -1384
rect 985 -1430 1145 -1417
rect 705 -1463 1145 -1430
rect 557 -1553 613 -1507
rect 705 -1553 1145 -1507
<< polycontact >>
rect -52 -1408 -6 -1361
rect 178 -1408 224 -1361
rect 865 -1430 985 -1384
<< metal1 >>
rect -169 -1450 -111 -1245
rect -52 -1361 -6 -1290
rect -52 -1420 -6 -1408
rect 178 -1361 224 -1290
rect 178 -1420 224 -1408
rect -179 -1465 -103 -1450
rect -179 -1512 -164 -1465
rect -118 -1512 -103 -1465
rect -179 -1527 -103 -1512
rect 48 -1465 124 -1450
rect 285 -1453 343 -1245
rect 742 -1384 1128 -1375
rect 742 -1430 865 -1384
rect 985 -1430 1128 -1384
rect 742 -1446 1128 -1430
rect 48 -1512 63 -1465
rect 109 -1512 124 -1465
rect 48 -1527 124 -1512
rect 275 -1468 351 -1453
rect 275 -1515 290 -1468
rect 336 -1515 351 -1468
rect 56 -1587 114 -1527
rect 275 -1530 351 -1515
rect 434 -1462 510 -1447
rect 434 -1509 449 -1462
rect 495 -1509 510 -1462
rect 434 -1524 510 -1509
rect 1193 -1462 1269 -1447
rect 1193 -1509 1208 -1462
rect 1254 -1509 1269 -1462
rect 1193 -1524 1269 -1509
rect 447 -1587 505 -1524
rect 56 -1634 505 -1587
rect 1201 -1690 1262 -1524
rect -229 -1805 1283 -1690
rect -229 -1806 76 -1805
<< labels >>
flabel metal1 -49 -1414 -9 -1307 1 FreeSans 400 0 0 0 INP
port 1 nsew signal input
flabel metal1 181 -1415 221 -1308 1 FreeSans 400 0 0 0 INN
port 2 nsew signal input
flabel metal1 -162 -1517 -118 -1261 1 FreeSans 400 0 0 0 OUTP
port 3 nsew power bidirectional
flabel metal1 291 -1524 335 -1268 1 FreeSans 400 0 0 0 OUTN
port 4 nsew power bidirectional
flabel metal1 766 -1433 1097 -1381 1 FreeSans 400 0 0 0 VBIAS
port 5 nsew power bidirectional
flabel metal1 1208 -1733 1255 -1458 1 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional
flabel pwell -219 -1801 19 -1695 1 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
<< end >>
